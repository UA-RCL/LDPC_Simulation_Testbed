CN_in_sig(344)	<=	VN_out_sig(0);
CN_in_sig(1512)	<=	VN_out_sig(1);
CN_in_sig(3816)	<=	VN_out_sig(2);
CN_in_sig(4872)	<=	VN_out_sig(3);
CN_in_sig(352)	<=	VN_out_sig(4);
CN_in_sig(1520)	<=	VN_out_sig(5);
CN_in_sig(3824)	<=	VN_out_sig(6);
CN_in_sig(4880)	<=	VN_out_sig(7);
CN_in_sig(360)	<=	VN_out_sig(8);
CN_in_sig(1528)	<=	VN_out_sig(9);
CN_in_sig(3832)	<=	VN_out_sig(10);
CN_in_sig(4888)	<=	VN_out_sig(11);
CN_in_sig(368)	<=	VN_out_sig(12);
CN_in_sig(1536)	<=	VN_out_sig(13);
CN_in_sig(3840)	<=	VN_out_sig(14);
CN_in_sig(4896)	<=	VN_out_sig(15);
CN_in_sig(376)	<=	VN_out_sig(16);
CN_in_sig(1544)	<=	VN_out_sig(17);
CN_in_sig(3848)	<=	VN_out_sig(18);
CN_in_sig(4904)	<=	VN_out_sig(19);
CN_in_sig(384)	<=	VN_out_sig(20);
CN_in_sig(1552)	<=	VN_out_sig(21);
CN_in_sig(3856)	<=	VN_out_sig(22);
CN_in_sig(4912)	<=	VN_out_sig(23);
CN_in_sig(392)	<=	VN_out_sig(24);
CN_in_sig(1560)	<=	VN_out_sig(25);
CN_in_sig(3864)	<=	VN_out_sig(26);
CN_in_sig(4920)	<=	VN_out_sig(27);
CN_in_sig(400)	<=	VN_out_sig(28);
CN_in_sig(1568)	<=	VN_out_sig(29);
CN_in_sig(3872)	<=	VN_out_sig(30);
CN_in_sig(4928)	<=	VN_out_sig(31);
CN_in_sig(408)	<=	VN_out_sig(32);
CN_in_sig(1576)	<=	VN_out_sig(33);
CN_in_sig(3880)	<=	VN_out_sig(34);
CN_in_sig(4936)	<=	VN_out_sig(35);
CN_in_sig(416)	<=	VN_out_sig(36);
CN_in_sig(1584)	<=	VN_out_sig(37);
CN_in_sig(3456)	<=	VN_out_sig(38);
CN_in_sig(4944)	<=	VN_out_sig(39);
CN_in_sig(424)	<=	VN_out_sig(40);
CN_in_sig(1592)	<=	VN_out_sig(41);
CN_in_sig(3464)	<=	VN_out_sig(42);
CN_in_sig(4952)	<=	VN_out_sig(43);
CN_in_sig(0)	<=	VN_out_sig(44);
CN_in_sig(1600)	<=	VN_out_sig(45);
CN_in_sig(3472)	<=	VN_out_sig(46);
CN_in_sig(4960)	<=	VN_out_sig(47);
CN_in_sig(8)	<=	VN_out_sig(48);
CN_in_sig(1608)	<=	VN_out_sig(49);
CN_in_sig(3480)	<=	VN_out_sig(50);
CN_in_sig(4968)	<=	VN_out_sig(51);
CN_in_sig(16)	<=	VN_out_sig(52);
CN_in_sig(1616)	<=	VN_out_sig(53);
CN_in_sig(3488)	<=	VN_out_sig(54);
CN_in_sig(4976)	<=	VN_out_sig(55);
CN_in_sig(24)	<=	VN_out_sig(56);
CN_in_sig(1624)	<=	VN_out_sig(57);
CN_in_sig(3496)	<=	VN_out_sig(58);
CN_in_sig(4984)	<=	VN_out_sig(59);
CN_in_sig(32)	<=	VN_out_sig(60);
CN_in_sig(1632)	<=	VN_out_sig(61);
CN_in_sig(3504)	<=	VN_out_sig(62);
CN_in_sig(4992)	<=	VN_out_sig(63);
CN_in_sig(40)	<=	VN_out_sig(64);
CN_in_sig(1640)	<=	VN_out_sig(65);
CN_in_sig(3512)	<=	VN_out_sig(66);
CN_in_sig(5000)	<=	VN_out_sig(67);
CN_in_sig(48)	<=	VN_out_sig(68);
CN_in_sig(1648)	<=	VN_out_sig(69);
CN_in_sig(3520)	<=	VN_out_sig(70);
CN_in_sig(5008)	<=	VN_out_sig(71);
CN_in_sig(56)	<=	VN_out_sig(72);
CN_in_sig(1656)	<=	VN_out_sig(73);
CN_in_sig(3528)	<=	VN_out_sig(74);
CN_in_sig(5016)	<=	VN_out_sig(75);
CN_in_sig(64)	<=	VN_out_sig(76);
CN_in_sig(1664)	<=	VN_out_sig(77);
CN_in_sig(3536)	<=	VN_out_sig(78);
CN_in_sig(5024)	<=	VN_out_sig(79);
CN_in_sig(72)	<=	VN_out_sig(80);
CN_in_sig(1672)	<=	VN_out_sig(81);
CN_in_sig(3544)	<=	VN_out_sig(82);
CN_in_sig(5032)	<=	VN_out_sig(83);
CN_in_sig(80)	<=	VN_out_sig(84);
CN_in_sig(1680)	<=	VN_out_sig(85);
CN_in_sig(3552)	<=	VN_out_sig(86);
CN_in_sig(5040)	<=	VN_out_sig(87);
CN_in_sig(88)	<=	VN_out_sig(88);
CN_in_sig(1688)	<=	VN_out_sig(89);
CN_in_sig(3560)	<=	VN_out_sig(90);
CN_in_sig(5048)	<=	VN_out_sig(91);
CN_in_sig(96)	<=	VN_out_sig(92);
CN_in_sig(1696)	<=	VN_out_sig(93);
CN_in_sig(3568)	<=	VN_out_sig(94);
CN_in_sig(5056)	<=	VN_out_sig(95);
CN_in_sig(104)	<=	VN_out_sig(96);
CN_in_sig(1704)	<=	VN_out_sig(97);
CN_in_sig(3576)	<=	VN_out_sig(98);
CN_in_sig(5064)	<=	VN_out_sig(99);
CN_in_sig(112)	<=	VN_out_sig(100);
CN_in_sig(1712)	<=	VN_out_sig(101);
CN_in_sig(3584)	<=	VN_out_sig(102);
CN_in_sig(5072)	<=	VN_out_sig(103);
CN_in_sig(120)	<=	VN_out_sig(104);
CN_in_sig(1720)	<=	VN_out_sig(105);
CN_in_sig(3592)	<=	VN_out_sig(106);
CN_in_sig(5080)	<=	VN_out_sig(107);
CN_in_sig(128)	<=	VN_out_sig(108);
CN_in_sig(1296)	<=	VN_out_sig(109);
CN_in_sig(3600)	<=	VN_out_sig(110);
CN_in_sig(5088)	<=	VN_out_sig(111);
CN_in_sig(136)	<=	VN_out_sig(112);
CN_in_sig(1304)	<=	VN_out_sig(113);
CN_in_sig(3608)	<=	VN_out_sig(114);
CN_in_sig(5096)	<=	VN_out_sig(115);
CN_in_sig(144)	<=	VN_out_sig(116);
CN_in_sig(1312)	<=	VN_out_sig(117);
CN_in_sig(3616)	<=	VN_out_sig(118);
CN_in_sig(5104)	<=	VN_out_sig(119);
CN_in_sig(152)	<=	VN_out_sig(120);
CN_in_sig(1320)	<=	VN_out_sig(121);
CN_in_sig(3624)	<=	VN_out_sig(122);
CN_in_sig(5112)	<=	VN_out_sig(123);
CN_in_sig(160)	<=	VN_out_sig(124);
CN_in_sig(1328)	<=	VN_out_sig(125);
CN_in_sig(3632)	<=	VN_out_sig(126);
CN_in_sig(5120)	<=	VN_out_sig(127);
CN_in_sig(168)	<=	VN_out_sig(128);
CN_in_sig(1336)	<=	VN_out_sig(129);
CN_in_sig(3640)	<=	VN_out_sig(130);
CN_in_sig(5128)	<=	VN_out_sig(131);
CN_in_sig(176)	<=	VN_out_sig(132);
CN_in_sig(1344)	<=	VN_out_sig(133);
CN_in_sig(3648)	<=	VN_out_sig(134);
CN_in_sig(5136)	<=	VN_out_sig(135);
CN_in_sig(184)	<=	VN_out_sig(136);
CN_in_sig(1352)	<=	VN_out_sig(137);
CN_in_sig(3656)	<=	VN_out_sig(138);
CN_in_sig(5144)	<=	VN_out_sig(139);
CN_in_sig(192)	<=	VN_out_sig(140);
CN_in_sig(1360)	<=	VN_out_sig(141);
CN_in_sig(3664)	<=	VN_out_sig(142);
CN_in_sig(5152)	<=	VN_out_sig(143);
CN_in_sig(200)	<=	VN_out_sig(144);
CN_in_sig(1368)	<=	VN_out_sig(145);
CN_in_sig(3672)	<=	VN_out_sig(146);
CN_in_sig(5160)	<=	VN_out_sig(147);
CN_in_sig(208)	<=	VN_out_sig(148);
CN_in_sig(1376)	<=	VN_out_sig(149);
CN_in_sig(3680)	<=	VN_out_sig(150);
CN_in_sig(5168)	<=	VN_out_sig(151);
CN_in_sig(216)	<=	VN_out_sig(152);
CN_in_sig(1384)	<=	VN_out_sig(153);
CN_in_sig(3688)	<=	VN_out_sig(154);
CN_in_sig(5176)	<=	VN_out_sig(155);
CN_in_sig(224)	<=	VN_out_sig(156);
CN_in_sig(1392)	<=	VN_out_sig(157);
CN_in_sig(3696)	<=	VN_out_sig(158);
CN_in_sig(4752)	<=	VN_out_sig(159);
CN_in_sig(232)	<=	VN_out_sig(160);
CN_in_sig(1400)	<=	VN_out_sig(161);
CN_in_sig(3704)	<=	VN_out_sig(162);
CN_in_sig(4760)	<=	VN_out_sig(163);
CN_in_sig(240)	<=	VN_out_sig(164);
CN_in_sig(1408)	<=	VN_out_sig(165);
CN_in_sig(3712)	<=	VN_out_sig(166);
CN_in_sig(4768)	<=	VN_out_sig(167);
CN_in_sig(248)	<=	VN_out_sig(168);
CN_in_sig(1416)	<=	VN_out_sig(169);
CN_in_sig(3720)	<=	VN_out_sig(170);
CN_in_sig(4776)	<=	VN_out_sig(171);
CN_in_sig(256)	<=	VN_out_sig(172);
CN_in_sig(1424)	<=	VN_out_sig(173);
CN_in_sig(3728)	<=	VN_out_sig(174);
CN_in_sig(4784)	<=	VN_out_sig(175);
CN_in_sig(264)	<=	VN_out_sig(176);
CN_in_sig(1432)	<=	VN_out_sig(177);
CN_in_sig(3736)	<=	VN_out_sig(178);
CN_in_sig(4792)	<=	VN_out_sig(179);
CN_in_sig(272)	<=	VN_out_sig(180);
CN_in_sig(1440)	<=	VN_out_sig(181);
CN_in_sig(3744)	<=	VN_out_sig(182);
CN_in_sig(4800)	<=	VN_out_sig(183);
CN_in_sig(280)	<=	VN_out_sig(184);
CN_in_sig(1448)	<=	VN_out_sig(185);
CN_in_sig(3752)	<=	VN_out_sig(186);
CN_in_sig(4808)	<=	VN_out_sig(187);
CN_in_sig(288)	<=	VN_out_sig(188);
CN_in_sig(1456)	<=	VN_out_sig(189);
CN_in_sig(3760)	<=	VN_out_sig(190);
CN_in_sig(4816)	<=	VN_out_sig(191);
CN_in_sig(296)	<=	VN_out_sig(192);
CN_in_sig(1464)	<=	VN_out_sig(193);
CN_in_sig(3768)	<=	VN_out_sig(194);
CN_in_sig(4824)	<=	VN_out_sig(195);
CN_in_sig(304)	<=	VN_out_sig(196);
CN_in_sig(1472)	<=	VN_out_sig(197);
CN_in_sig(3776)	<=	VN_out_sig(198);
CN_in_sig(4832)	<=	VN_out_sig(199);
CN_in_sig(312)	<=	VN_out_sig(200);
CN_in_sig(1480)	<=	VN_out_sig(201);
CN_in_sig(3784)	<=	VN_out_sig(202);
CN_in_sig(4840)	<=	VN_out_sig(203);
CN_in_sig(320)	<=	VN_out_sig(204);
CN_in_sig(1488)	<=	VN_out_sig(205);
CN_in_sig(3792)	<=	VN_out_sig(206);
CN_in_sig(4848)	<=	VN_out_sig(207);
CN_in_sig(328)	<=	VN_out_sig(208);
CN_in_sig(1496)	<=	VN_out_sig(209);
CN_in_sig(3800)	<=	VN_out_sig(210);
CN_in_sig(4856)	<=	VN_out_sig(211);
CN_in_sig(336)	<=	VN_out_sig(212);
CN_in_sig(1504)	<=	VN_out_sig(213);
CN_in_sig(3808)	<=	VN_out_sig(214);
CN_in_sig(4864)	<=	VN_out_sig(215);
CN_in_sig(664)	<=	VN_out_sig(216);
CN_in_sig(1824)	<=	VN_out_sig(217);
CN_in_sig(3224)	<=	VN_out_sig(218);
CN_in_sig(4720)	<=	VN_out_sig(219);
CN_in_sig(672)	<=	VN_out_sig(220);
CN_in_sig(1832)	<=	VN_out_sig(221);
CN_in_sig(3232)	<=	VN_out_sig(222);
CN_in_sig(4728)	<=	VN_out_sig(223);
CN_in_sig(680)	<=	VN_out_sig(224);
CN_in_sig(1840)	<=	VN_out_sig(225);
CN_in_sig(3240)	<=	VN_out_sig(226);
CN_in_sig(4736)	<=	VN_out_sig(227);
CN_in_sig(688)	<=	VN_out_sig(228);
CN_in_sig(1848)	<=	VN_out_sig(229);
CN_in_sig(3248)	<=	VN_out_sig(230);
CN_in_sig(4744)	<=	VN_out_sig(231);
CN_in_sig(696)	<=	VN_out_sig(232);
CN_in_sig(1856)	<=	VN_out_sig(233);
CN_in_sig(3256)	<=	VN_out_sig(234);
CN_in_sig(4320)	<=	VN_out_sig(235);
CN_in_sig(704)	<=	VN_out_sig(236);
CN_in_sig(1864)	<=	VN_out_sig(237);
CN_in_sig(3264)	<=	VN_out_sig(238);
CN_in_sig(4328)	<=	VN_out_sig(239);
CN_in_sig(712)	<=	VN_out_sig(240);
CN_in_sig(1872)	<=	VN_out_sig(241);
CN_in_sig(3272)	<=	VN_out_sig(242);
CN_in_sig(4336)	<=	VN_out_sig(243);
CN_in_sig(720)	<=	VN_out_sig(244);
CN_in_sig(1880)	<=	VN_out_sig(245);
CN_in_sig(3280)	<=	VN_out_sig(246);
CN_in_sig(4344)	<=	VN_out_sig(247);
CN_in_sig(728)	<=	VN_out_sig(248);
CN_in_sig(1888)	<=	VN_out_sig(249);
CN_in_sig(3288)	<=	VN_out_sig(250);
CN_in_sig(4352)	<=	VN_out_sig(251);
CN_in_sig(736)	<=	VN_out_sig(252);
CN_in_sig(1896)	<=	VN_out_sig(253);
CN_in_sig(3296)	<=	VN_out_sig(254);
CN_in_sig(4360)	<=	VN_out_sig(255);
CN_in_sig(744)	<=	VN_out_sig(256);
CN_in_sig(1904)	<=	VN_out_sig(257);
CN_in_sig(3304)	<=	VN_out_sig(258);
CN_in_sig(4368)	<=	VN_out_sig(259);
CN_in_sig(752)	<=	VN_out_sig(260);
CN_in_sig(1912)	<=	VN_out_sig(261);
CN_in_sig(3312)	<=	VN_out_sig(262);
CN_in_sig(4376)	<=	VN_out_sig(263);
CN_in_sig(760)	<=	VN_out_sig(264);
CN_in_sig(1920)	<=	VN_out_sig(265);
CN_in_sig(3320)	<=	VN_out_sig(266);
CN_in_sig(4384)	<=	VN_out_sig(267);
CN_in_sig(768)	<=	VN_out_sig(268);
CN_in_sig(1928)	<=	VN_out_sig(269);
CN_in_sig(3328)	<=	VN_out_sig(270);
CN_in_sig(4392)	<=	VN_out_sig(271);
CN_in_sig(776)	<=	VN_out_sig(272);
CN_in_sig(1936)	<=	VN_out_sig(273);
CN_in_sig(3336)	<=	VN_out_sig(274);
CN_in_sig(4400)	<=	VN_out_sig(275);
CN_in_sig(784)	<=	VN_out_sig(276);
CN_in_sig(1944)	<=	VN_out_sig(277);
CN_in_sig(3344)	<=	VN_out_sig(278);
CN_in_sig(4408)	<=	VN_out_sig(279);
CN_in_sig(792)	<=	VN_out_sig(280);
CN_in_sig(1952)	<=	VN_out_sig(281);
CN_in_sig(3352)	<=	VN_out_sig(282);
CN_in_sig(4416)	<=	VN_out_sig(283);
CN_in_sig(800)	<=	VN_out_sig(284);
CN_in_sig(1960)	<=	VN_out_sig(285);
CN_in_sig(3360)	<=	VN_out_sig(286);
CN_in_sig(4424)	<=	VN_out_sig(287);
CN_in_sig(808)	<=	VN_out_sig(288);
CN_in_sig(1968)	<=	VN_out_sig(289);
CN_in_sig(3368)	<=	VN_out_sig(290);
CN_in_sig(4432)	<=	VN_out_sig(291);
CN_in_sig(816)	<=	VN_out_sig(292);
CN_in_sig(1976)	<=	VN_out_sig(293);
CN_in_sig(3376)	<=	VN_out_sig(294);
CN_in_sig(4440)	<=	VN_out_sig(295);
CN_in_sig(824)	<=	VN_out_sig(296);
CN_in_sig(1984)	<=	VN_out_sig(297);
CN_in_sig(3384)	<=	VN_out_sig(298);
CN_in_sig(4448)	<=	VN_out_sig(299);
CN_in_sig(832)	<=	VN_out_sig(300);
CN_in_sig(1992)	<=	VN_out_sig(301);
CN_in_sig(3392)	<=	VN_out_sig(302);
CN_in_sig(4456)	<=	VN_out_sig(303);
CN_in_sig(840)	<=	VN_out_sig(304);
CN_in_sig(2000)	<=	VN_out_sig(305);
CN_in_sig(3400)	<=	VN_out_sig(306);
CN_in_sig(4464)	<=	VN_out_sig(307);
CN_in_sig(848)	<=	VN_out_sig(308);
CN_in_sig(2008)	<=	VN_out_sig(309);
CN_in_sig(3408)	<=	VN_out_sig(310);
CN_in_sig(4472)	<=	VN_out_sig(311);
CN_in_sig(856)	<=	VN_out_sig(312);
CN_in_sig(2016)	<=	VN_out_sig(313);
CN_in_sig(3416)	<=	VN_out_sig(314);
CN_in_sig(4480)	<=	VN_out_sig(315);
CN_in_sig(432)	<=	VN_out_sig(316);
CN_in_sig(2024)	<=	VN_out_sig(317);
CN_in_sig(3424)	<=	VN_out_sig(318);
CN_in_sig(4488)	<=	VN_out_sig(319);
CN_in_sig(440)	<=	VN_out_sig(320);
CN_in_sig(2032)	<=	VN_out_sig(321);
CN_in_sig(3432)	<=	VN_out_sig(322);
CN_in_sig(4496)	<=	VN_out_sig(323);
CN_in_sig(448)	<=	VN_out_sig(324);
CN_in_sig(2040)	<=	VN_out_sig(325);
CN_in_sig(3440)	<=	VN_out_sig(326);
CN_in_sig(4504)	<=	VN_out_sig(327);
CN_in_sig(456)	<=	VN_out_sig(328);
CN_in_sig(2048)	<=	VN_out_sig(329);
CN_in_sig(3448)	<=	VN_out_sig(330);
CN_in_sig(4512)	<=	VN_out_sig(331);
CN_in_sig(464)	<=	VN_out_sig(332);
CN_in_sig(2056)	<=	VN_out_sig(333);
CN_in_sig(3024)	<=	VN_out_sig(334);
CN_in_sig(4520)	<=	VN_out_sig(335);
CN_in_sig(472)	<=	VN_out_sig(336);
CN_in_sig(2064)	<=	VN_out_sig(337);
CN_in_sig(3032)	<=	VN_out_sig(338);
CN_in_sig(4528)	<=	VN_out_sig(339);
CN_in_sig(480)	<=	VN_out_sig(340);
CN_in_sig(2072)	<=	VN_out_sig(341);
CN_in_sig(3040)	<=	VN_out_sig(342);
CN_in_sig(4536)	<=	VN_out_sig(343);
CN_in_sig(488)	<=	VN_out_sig(344);
CN_in_sig(2080)	<=	VN_out_sig(345);
CN_in_sig(3048)	<=	VN_out_sig(346);
CN_in_sig(4544)	<=	VN_out_sig(347);
CN_in_sig(496)	<=	VN_out_sig(348);
CN_in_sig(2088)	<=	VN_out_sig(349);
CN_in_sig(3056)	<=	VN_out_sig(350);
CN_in_sig(4552)	<=	VN_out_sig(351);
CN_in_sig(504)	<=	VN_out_sig(352);
CN_in_sig(2096)	<=	VN_out_sig(353);
CN_in_sig(3064)	<=	VN_out_sig(354);
CN_in_sig(4560)	<=	VN_out_sig(355);
CN_in_sig(512)	<=	VN_out_sig(356);
CN_in_sig(2104)	<=	VN_out_sig(357);
CN_in_sig(3072)	<=	VN_out_sig(358);
CN_in_sig(4568)	<=	VN_out_sig(359);
CN_in_sig(520)	<=	VN_out_sig(360);
CN_in_sig(2112)	<=	VN_out_sig(361);
CN_in_sig(3080)	<=	VN_out_sig(362);
CN_in_sig(4576)	<=	VN_out_sig(363);
CN_in_sig(528)	<=	VN_out_sig(364);
CN_in_sig(2120)	<=	VN_out_sig(365);
CN_in_sig(3088)	<=	VN_out_sig(366);
CN_in_sig(4584)	<=	VN_out_sig(367);
CN_in_sig(536)	<=	VN_out_sig(368);
CN_in_sig(2128)	<=	VN_out_sig(369);
CN_in_sig(3096)	<=	VN_out_sig(370);
CN_in_sig(4592)	<=	VN_out_sig(371);
CN_in_sig(544)	<=	VN_out_sig(372);
CN_in_sig(2136)	<=	VN_out_sig(373);
CN_in_sig(3104)	<=	VN_out_sig(374);
CN_in_sig(4600)	<=	VN_out_sig(375);
CN_in_sig(552)	<=	VN_out_sig(376);
CN_in_sig(2144)	<=	VN_out_sig(377);
CN_in_sig(3112)	<=	VN_out_sig(378);
CN_in_sig(4608)	<=	VN_out_sig(379);
CN_in_sig(560)	<=	VN_out_sig(380);
CN_in_sig(2152)	<=	VN_out_sig(381);
CN_in_sig(3120)	<=	VN_out_sig(382);
CN_in_sig(4616)	<=	VN_out_sig(383);
CN_in_sig(568)	<=	VN_out_sig(384);
CN_in_sig(1728)	<=	VN_out_sig(385);
CN_in_sig(3128)	<=	VN_out_sig(386);
CN_in_sig(4624)	<=	VN_out_sig(387);
CN_in_sig(576)	<=	VN_out_sig(388);
CN_in_sig(1736)	<=	VN_out_sig(389);
CN_in_sig(3136)	<=	VN_out_sig(390);
CN_in_sig(4632)	<=	VN_out_sig(391);
CN_in_sig(584)	<=	VN_out_sig(392);
CN_in_sig(1744)	<=	VN_out_sig(393);
CN_in_sig(3144)	<=	VN_out_sig(394);
CN_in_sig(4640)	<=	VN_out_sig(395);
CN_in_sig(592)	<=	VN_out_sig(396);
CN_in_sig(1752)	<=	VN_out_sig(397);
CN_in_sig(3152)	<=	VN_out_sig(398);
CN_in_sig(4648)	<=	VN_out_sig(399);
CN_in_sig(600)	<=	VN_out_sig(400);
CN_in_sig(1760)	<=	VN_out_sig(401);
CN_in_sig(3160)	<=	VN_out_sig(402);
CN_in_sig(4656)	<=	VN_out_sig(403);
CN_in_sig(608)	<=	VN_out_sig(404);
CN_in_sig(1768)	<=	VN_out_sig(405);
CN_in_sig(3168)	<=	VN_out_sig(406);
CN_in_sig(4664)	<=	VN_out_sig(407);
CN_in_sig(616)	<=	VN_out_sig(408);
CN_in_sig(1776)	<=	VN_out_sig(409);
CN_in_sig(3176)	<=	VN_out_sig(410);
CN_in_sig(4672)	<=	VN_out_sig(411);
CN_in_sig(624)	<=	VN_out_sig(412);
CN_in_sig(1784)	<=	VN_out_sig(413);
CN_in_sig(3184)	<=	VN_out_sig(414);
CN_in_sig(4680)	<=	VN_out_sig(415);
CN_in_sig(632)	<=	VN_out_sig(416);
CN_in_sig(1792)	<=	VN_out_sig(417);
CN_in_sig(3192)	<=	VN_out_sig(418);
CN_in_sig(4688)	<=	VN_out_sig(419);
CN_in_sig(640)	<=	VN_out_sig(420);
CN_in_sig(1800)	<=	VN_out_sig(421);
CN_in_sig(3200)	<=	VN_out_sig(422);
CN_in_sig(4696)	<=	VN_out_sig(423);
CN_in_sig(648)	<=	VN_out_sig(424);
CN_in_sig(1808)	<=	VN_out_sig(425);
CN_in_sig(3208)	<=	VN_out_sig(426);
CN_in_sig(4704)	<=	VN_out_sig(427);
CN_in_sig(656)	<=	VN_out_sig(428);
CN_in_sig(1816)	<=	VN_out_sig(429);
CN_in_sig(3216)	<=	VN_out_sig(430);
CN_in_sig(4712)	<=	VN_out_sig(431);
CN_in_sig(944)	<=	VN_out_sig(432);
CN_in_sig(2400)	<=	VN_out_sig(433);
CN_in_sig(2704)	<=	VN_out_sig(434);
CN_in_sig(3896)	<=	VN_out_sig(435);
CN_in_sig(952)	<=	VN_out_sig(436);
CN_in_sig(2408)	<=	VN_out_sig(437);
CN_in_sig(2712)	<=	VN_out_sig(438);
CN_in_sig(3904)	<=	VN_out_sig(439);
CN_in_sig(960)	<=	VN_out_sig(440);
CN_in_sig(2416)	<=	VN_out_sig(441);
CN_in_sig(2720)	<=	VN_out_sig(442);
CN_in_sig(3912)	<=	VN_out_sig(443);
CN_in_sig(968)	<=	VN_out_sig(444);
CN_in_sig(2424)	<=	VN_out_sig(445);
CN_in_sig(2728)	<=	VN_out_sig(446);
CN_in_sig(3920)	<=	VN_out_sig(447);
CN_in_sig(976)	<=	VN_out_sig(448);
CN_in_sig(2432)	<=	VN_out_sig(449);
CN_in_sig(2736)	<=	VN_out_sig(450);
CN_in_sig(3928)	<=	VN_out_sig(451);
CN_in_sig(984)	<=	VN_out_sig(452);
CN_in_sig(2440)	<=	VN_out_sig(453);
CN_in_sig(2744)	<=	VN_out_sig(454);
CN_in_sig(3936)	<=	VN_out_sig(455);
CN_in_sig(992)	<=	VN_out_sig(456);
CN_in_sig(2448)	<=	VN_out_sig(457);
CN_in_sig(2752)	<=	VN_out_sig(458);
CN_in_sig(3944)	<=	VN_out_sig(459);
CN_in_sig(1000)	<=	VN_out_sig(460);
CN_in_sig(2456)	<=	VN_out_sig(461);
CN_in_sig(2760)	<=	VN_out_sig(462);
CN_in_sig(3952)	<=	VN_out_sig(463);
CN_in_sig(1008)	<=	VN_out_sig(464);
CN_in_sig(2464)	<=	VN_out_sig(465);
CN_in_sig(2768)	<=	VN_out_sig(466);
CN_in_sig(3960)	<=	VN_out_sig(467);
CN_in_sig(1016)	<=	VN_out_sig(468);
CN_in_sig(2472)	<=	VN_out_sig(469);
CN_in_sig(2776)	<=	VN_out_sig(470);
CN_in_sig(3968)	<=	VN_out_sig(471);
CN_in_sig(1024)	<=	VN_out_sig(472);
CN_in_sig(2480)	<=	VN_out_sig(473);
CN_in_sig(2784)	<=	VN_out_sig(474);
CN_in_sig(3976)	<=	VN_out_sig(475);
CN_in_sig(1032)	<=	VN_out_sig(476);
CN_in_sig(2488)	<=	VN_out_sig(477);
CN_in_sig(2792)	<=	VN_out_sig(478);
CN_in_sig(3984)	<=	VN_out_sig(479);
CN_in_sig(1040)	<=	VN_out_sig(480);
CN_in_sig(2496)	<=	VN_out_sig(481);
CN_in_sig(2800)	<=	VN_out_sig(482);
CN_in_sig(3992)	<=	VN_out_sig(483);
CN_in_sig(1048)	<=	VN_out_sig(484);
CN_in_sig(2504)	<=	VN_out_sig(485);
CN_in_sig(2808)	<=	VN_out_sig(486);
CN_in_sig(4000)	<=	VN_out_sig(487);
CN_in_sig(1056)	<=	VN_out_sig(488);
CN_in_sig(2512)	<=	VN_out_sig(489);
CN_in_sig(2816)	<=	VN_out_sig(490);
CN_in_sig(4008)	<=	VN_out_sig(491);
CN_in_sig(1064)	<=	VN_out_sig(492);
CN_in_sig(2520)	<=	VN_out_sig(493);
CN_in_sig(2824)	<=	VN_out_sig(494);
CN_in_sig(4016)	<=	VN_out_sig(495);
CN_in_sig(1072)	<=	VN_out_sig(496);
CN_in_sig(2528)	<=	VN_out_sig(497);
CN_in_sig(2832)	<=	VN_out_sig(498);
CN_in_sig(4024)	<=	VN_out_sig(499);
CN_in_sig(1080)	<=	VN_out_sig(500);
CN_in_sig(2536)	<=	VN_out_sig(501);
CN_in_sig(2840)	<=	VN_out_sig(502);
CN_in_sig(4032)	<=	VN_out_sig(503);
CN_in_sig(1088)	<=	VN_out_sig(504);
CN_in_sig(2544)	<=	VN_out_sig(505);
CN_in_sig(2848)	<=	VN_out_sig(506);
CN_in_sig(4040)	<=	VN_out_sig(507);
CN_in_sig(1096)	<=	VN_out_sig(508);
CN_in_sig(2552)	<=	VN_out_sig(509);
CN_in_sig(2856)	<=	VN_out_sig(510);
CN_in_sig(4048)	<=	VN_out_sig(511);
CN_in_sig(1104)	<=	VN_out_sig(512);
CN_in_sig(2560)	<=	VN_out_sig(513);
CN_in_sig(2864)	<=	VN_out_sig(514);
CN_in_sig(4056)	<=	VN_out_sig(515);
CN_in_sig(1112)	<=	VN_out_sig(516);
CN_in_sig(2568)	<=	VN_out_sig(517);
CN_in_sig(2872)	<=	VN_out_sig(518);
CN_in_sig(4064)	<=	VN_out_sig(519);
CN_in_sig(1120)	<=	VN_out_sig(520);
CN_in_sig(2576)	<=	VN_out_sig(521);
CN_in_sig(2880)	<=	VN_out_sig(522);
CN_in_sig(4072)	<=	VN_out_sig(523);
CN_in_sig(1128)	<=	VN_out_sig(524);
CN_in_sig(2584)	<=	VN_out_sig(525);
CN_in_sig(2888)	<=	VN_out_sig(526);
CN_in_sig(4080)	<=	VN_out_sig(527);
CN_in_sig(1136)	<=	VN_out_sig(528);
CN_in_sig(2160)	<=	VN_out_sig(529);
CN_in_sig(2896)	<=	VN_out_sig(530);
CN_in_sig(4088)	<=	VN_out_sig(531);
CN_in_sig(1144)	<=	VN_out_sig(532);
CN_in_sig(2168)	<=	VN_out_sig(533);
CN_in_sig(2904)	<=	VN_out_sig(534);
CN_in_sig(4096)	<=	VN_out_sig(535);
CN_in_sig(1152)	<=	VN_out_sig(536);
CN_in_sig(2176)	<=	VN_out_sig(537);
CN_in_sig(2912)	<=	VN_out_sig(538);
CN_in_sig(4104)	<=	VN_out_sig(539);
CN_in_sig(1160)	<=	VN_out_sig(540);
CN_in_sig(2184)	<=	VN_out_sig(541);
CN_in_sig(2920)	<=	VN_out_sig(542);
CN_in_sig(4112)	<=	VN_out_sig(543);
CN_in_sig(1168)	<=	VN_out_sig(544);
CN_in_sig(2192)	<=	VN_out_sig(545);
CN_in_sig(2928)	<=	VN_out_sig(546);
CN_in_sig(4120)	<=	VN_out_sig(547);
CN_in_sig(1176)	<=	VN_out_sig(548);
CN_in_sig(2200)	<=	VN_out_sig(549);
CN_in_sig(2936)	<=	VN_out_sig(550);
CN_in_sig(4128)	<=	VN_out_sig(551);
CN_in_sig(1184)	<=	VN_out_sig(552);
CN_in_sig(2208)	<=	VN_out_sig(553);
CN_in_sig(2944)	<=	VN_out_sig(554);
CN_in_sig(4136)	<=	VN_out_sig(555);
CN_in_sig(1192)	<=	VN_out_sig(556);
CN_in_sig(2216)	<=	VN_out_sig(557);
CN_in_sig(2952)	<=	VN_out_sig(558);
CN_in_sig(4144)	<=	VN_out_sig(559);
CN_in_sig(1200)	<=	VN_out_sig(560);
CN_in_sig(2224)	<=	VN_out_sig(561);
CN_in_sig(2960)	<=	VN_out_sig(562);
CN_in_sig(4152)	<=	VN_out_sig(563);
CN_in_sig(1208)	<=	VN_out_sig(564);
CN_in_sig(2232)	<=	VN_out_sig(565);
CN_in_sig(2968)	<=	VN_out_sig(566);
CN_in_sig(4160)	<=	VN_out_sig(567);
CN_in_sig(1216)	<=	VN_out_sig(568);
CN_in_sig(2240)	<=	VN_out_sig(569);
CN_in_sig(2976)	<=	VN_out_sig(570);
CN_in_sig(4168)	<=	VN_out_sig(571);
CN_in_sig(1224)	<=	VN_out_sig(572);
CN_in_sig(2248)	<=	VN_out_sig(573);
CN_in_sig(2984)	<=	VN_out_sig(574);
CN_in_sig(4176)	<=	VN_out_sig(575);
CN_in_sig(1232)	<=	VN_out_sig(576);
CN_in_sig(2256)	<=	VN_out_sig(577);
CN_in_sig(2992)	<=	VN_out_sig(578);
CN_in_sig(4184)	<=	VN_out_sig(579);
CN_in_sig(1240)	<=	VN_out_sig(580);
CN_in_sig(2264)	<=	VN_out_sig(581);
CN_in_sig(3000)	<=	VN_out_sig(582);
CN_in_sig(4192)	<=	VN_out_sig(583);
CN_in_sig(1248)	<=	VN_out_sig(584);
CN_in_sig(2272)	<=	VN_out_sig(585);
CN_in_sig(3008)	<=	VN_out_sig(586);
CN_in_sig(4200)	<=	VN_out_sig(587);
CN_in_sig(1256)	<=	VN_out_sig(588);
CN_in_sig(2280)	<=	VN_out_sig(589);
CN_in_sig(3016)	<=	VN_out_sig(590);
CN_in_sig(4208)	<=	VN_out_sig(591);
CN_in_sig(1264)	<=	VN_out_sig(592);
CN_in_sig(2288)	<=	VN_out_sig(593);
CN_in_sig(2592)	<=	VN_out_sig(594);
CN_in_sig(4216)	<=	VN_out_sig(595);
CN_in_sig(1272)	<=	VN_out_sig(596);
CN_in_sig(2296)	<=	VN_out_sig(597);
CN_in_sig(2600)	<=	VN_out_sig(598);
CN_in_sig(4224)	<=	VN_out_sig(599);
CN_in_sig(1280)	<=	VN_out_sig(600);
CN_in_sig(2304)	<=	VN_out_sig(601);
CN_in_sig(2608)	<=	VN_out_sig(602);
CN_in_sig(4232)	<=	VN_out_sig(603);
CN_in_sig(1288)	<=	VN_out_sig(604);
CN_in_sig(2312)	<=	VN_out_sig(605);
CN_in_sig(2616)	<=	VN_out_sig(606);
CN_in_sig(4240)	<=	VN_out_sig(607);
CN_in_sig(864)	<=	VN_out_sig(608);
CN_in_sig(2320)	<=	VN_out_sig(609);
CN_in_sig(2624)	<=	VN_out_sig(610);
CN_in_sig(4248)	<=	VN_out_sig(611);
CN_in_sig(872)	<=	VN_out_sig(612);
CN_in_sig(2328)	<=	VN_out_sig(613);
CN_in_sig(2632)	<=	VN_out_sig(614);
CN_in_sig(4256)	<=	VN_out_sig(615);
CN_in_sig(880)	<=	VN_out_sig(616);
CN_in_sig(2336)	<=	VN_out_sig(617);
CN_in_sig(2640)	<=	VN_out_sig(618);
CN_in_sig(4264)	<=	VN_out_sig(619);
CN_in_sig(888)	<=	VN_out_sig(620);
CN_in_sig(2344)	<=	VN_out_sig(621);
CN_in_sig(2648)	<=	VN_out_sig(622);
CN_in_sig(4272)	<=	VN_out_sig(623);
CN_in_sig(896)	<=	VN_out_sig(624);
CN_in_sig(2352)	<=	VN_out_sig(625);
CN_in_sig(2656)	<=	VN_out_sig(626);
CN_in_sig(4280)	<=	VN_out_sig(627);
CN_in_sig(904)	<=	VN_out_sig(628);
CN_in_sig(2360)	<=	VN_out_sig(629);
CN_in_sig(2664)	<=	VN_out_sig(630);
CN_in_sig(4288)	<=	VN_out_sig(631);
CN_in_sig(912)	<=	VN_out_sig(632);
CN_in_sig(2368)	<=	VN_out_sig(633);
CN_in_sig(2672)	<=	VN_out_sig(634);
CN_in_sig(4296)	<=	VN_out_sig(635);
CN_in_sig(920)	<=	VN_out_sig(636);
CN_in_sig(2376)	<=	VN_out_sig(637);
CN_in_sig(2680)	<=	VN_out_sig(638);
CN_in_sig(4304)	<=	VN_out_sig(639);
CN_in_sig(928)	<=	VN_out_sig(640);
CN_in_sig(2384)	<=	VN_out_sig(641);
CN_in_sig(2688)	<=	VN_out_sig(642);
CN_in_sig(4312)	<=	VN_out_sig(643);
CN_in_sig(936)	<=	VN_out_sig(644);
CN_in_sig(2392)	<=	VN_out_sig(645);
CN_in_sig(2696)	<=	VN_out_sig(646);
CN_in_sig(3888)	<=	VN_out_sig(647);
CN_in_sig(1265)	<=	VN_out_sig(648);
CN_in_sig(1985)	<=	VN_out_sig(649);
CN_in_sig(3025)	<=	VN_out_sig(650);
CN_in_sig(5049)	<=	VN_out_sig(651);
CN_in_sig(1273)	<=	VN_out_sig(652);
CN_in_sig(1993)	<=	VN_out_sig(653);
CN_in_sig(3033)	<=	VN_out_sig(654);
CN_in_sig(5057)	<=	VN_out_sig(655);
CN_in_sig(1281)	<=	VN_out_sig(656);
CN_in_sig(2001)	<=	VN_out_sig(657);
CN_in_sig(3041)	<=	VN_out_sig(658);
CN_in_sig(5065)	<=	VN_out_sig(659);
CN_in_sig(1289)	<=	VN_out_sig(660);
CN_in_sig(2009)	<=	VN_out_sig(661);
CN_in_sig(3049)	<=	VN_out_sig(662);
CN_in_sig(5073)	<=	VN_out_sig(663);
CN_in_sig(865)	<=	VN_out_sig(664);
CN_in_sig(2017)	<=	VN_out_sig(665);
CN_in_sig(3057)	<=	VN_out_sig(666);
CN_in_sig(5081)	<=	VN_out_sig(667);
CN_in_sig(873)	<=	VN_out_sig(668);
CN_in_sig(2025)	<=	VN_out_sig(669);
CN_in_sig(3065)	<=	VN_out_sig(670);
CN_in_sig(5089)	<=	VN_out_sig(671);
CN_in_sig(881)	<=	VN_out_sig(672);
CN_in_sig(2033)	<=	VN_out_sig(673);
CN_in_sig(3073)	<=	VN_out_sig(674);
CN_in_sig(5097)	<=	VN_out_sig(675);
CN_in_sig(889)	<=	VN_out_sig(676);
CN_in_sig(2041)	<=	VN_out_sig(677);
CN_in_sig(3081)	<=	VN_out_sig(678);
CN_in_sig(5105)	<=	VN_out_sig(679);
CN_in_sig(897)	<=	VN_out_sig(680);
CN_in_sig(2049)	<=	VN_out_sig(681);
CN_in_sig(3089)	<=	VN_out_sig(682);
CN_in_sig(5113)	<=	VN_out_sig(683);
CN_in_sig(905)	<=	VN_out_sig(684);
CN_in_sig(2057)	<=	VN_out_sig(685);
CN_in_sig(3097)	<=	VN_out_sig(686);
CN_in_sig(5121)	<=	VN_out_sig(687);
CN_in_sig(913)	<=	VN_out_sig(688);
CN_in_sig(2065)	<=	VN_out_sig(689);
CN_in_sig(3105)	<=	VN_out_sig(690);
CN_in_sig(5129)	<=	VN_out_sig(691);
CN_in_sig(921)	<=	VN_out_sig(692);
CN_in_sig(2073)	<=	VN_out_sig(693);
CN_in_sig(3113)	<=	VN_out_sig(694);
CN_in_sig(5137)	<=	VN_out_sig(695);
CN_in_sig(929)	<=	VN_out_sig(696);
CN_in_sig(2081)	<=	VN_out_sig(697);
CN_in_sig(3121)	<=	VN_out_sig(698);
CN_in_sig(5145)	<=	VN_out_sig(699);
CN_in_sig(937)	<=	VN_out_sig(700);
CN_in_sig(2089)	<=	VN_out_sig(701);
CN_in_sig(3129)	<=	VN_out_sig(702);
CN_in_sig(5153)	<=	VN_out_sig(703);
CN_in_sig(945)	<=	VN_out_sig(704);
CN_in_sig(2097)	<=	VN_out_sig(705);
CN_in_sig(3137)	<=	VN_out_sig(706);
CN_in_sig(5161)	<=	VN_out_sig(707);
CN_in_sig(953)	<=	VN_out_sig(708);
CN_in_sig(2105)	<=	VN_out_sig(709);
CN_in_sig(3145)	<=	VN_out_sig(710);
CN_in_sig(5169)	<=	VN_out_sig(711);
CN_in_sig(961)	<=	VN_out_sig(712);
CN_in_sig(2113)	<=	VN_out_sig(713);
CN_in_sig(3153)	<=	VN_out_sig(714);
CN_in_sig(5177)	<=	VN_out_sig(715);
CN_in_sig(969)	<=	VN_out_sig(716);
CN_in_sig(2121)	<=	VN_out_sig(717);
CN_in_sig(3161)	<=	VN_out_sig(718);
CN_in_sig(4753)	<=	VN_out_sig(719);
CN_in_sig(977)	<=	VN_out_sig(720);
CN_in_sig(2129)	<=	VN_out_sig(721);
CN_in_sig(3169)	<=	VN_out_sig(722);
CN_in_sig(4761)	<=	VN_out_sig(723);
CN_in_sig(985)	<=	VN_out_sig(724);
CN_in_sig(2137)	<=	VN_out_sig(725);
CN_in_sig(3177)	<=	VN_out_sig(726);
CN_in_sig(4769)	<=	VN_out_sig(727);
CN_in_sig(993)	<=	VN_out_sig(728);
CN_in_sig(2145)	<=	VN_out_sig(729);
CN_in_sig(3185)	<=	VN_out_sig(730);
CN_in_sig(4777)	<=	VN_out_sig(731);
CN_in_sig(1001)	<=	VN_out_sig(732);
CN_in_sig(2153)	<=	VN_out_sig(733);
CN_in_sig(3193)	<=	VN_out_sig(734);
CN_in_sig(4785)	<=	VN_out_sig(735);
CN_in_sig(1009)	<=	VN_out_sig(736);
CN_in_sig(1729)	<=	VN_out_sig(737);
CN_in_sig(3201)	<=	VN_out_sig(738);
CN_in_sig(4793)	<=	VN_out_sig(739);
CN_in_sig(1017)	<=	VN_out_sig(740);
CN_in_sig(1737)	<=	VN_out_sig(741);
CN_in_sig(3209)	<=	VN_out_sig(742);
CN_in_sig(4801)	<=	VN_out_sig(743);
CN_in_sig(1025)	<=	VN_out_sig(744);
CN_in_sig(1745)	<=	VN_out_sig(745);
CN_in_sig(3217)	<=	VN_out_sig(746);
CN_in_sig(4809)	<=	VN_out_sig(747);
CN_in_sig(1033)	<=	VN_out_sig(748);
CN_in_sig(1753)	<=	VN_out_sig(749);
CN_in_sig(3225)	<=	VN_out_sig(750);
CN_in_sig(4817)	<=	VN_out_sig(751);
CN_in_sig(1041)	<=	VN_out_sig(752);
CN_in_sig(1761)	<=	VN_out_sig(753);
CN_in_sig(3233)	<=	VN_out_sig(754);
CN_in_sig(4825)	<=	VN_out_sig(755);
CN_in_sig(1049)	<=	VN_out_sig(756);
CN_in_sig(1769)	<=	VN_out_sig(757);
CN_in_sig(3241)	<=	VN_out_sig(758);
CN_in_sig(4833)	<=	VN_out_sig(759);
CN_in_sig(1057)	<=	VN_out_sig(760);
CN_in_sig(1777)	<=	VN_out_sig(761);
CN_in_sig(3249)	<=	VN_out_sig(762);
CN_in_sig(4841)	<=	VN_out_sig(763);
CN_in_sig(1065)	<=	VN_out_sig(764);
CN_in_sig(1785)	<=	VN_out_sig(765);
CN_in_sig(3257)	<=	VN_out_sig(766);
CN_in_sig(4849)	<=	VN_out_sig(767);
CN_in_sig(1073)	<=	VN_out_sig(768);
CN_in_sig(1793)	<=	VN_out_sig(769);
CN_in_sig(3265)	<=	VN_out_sig(770);
CN_in_sig(4857)	<=	VN_out_sig(771);
CN_in_sig(1081)	<=	VN_out_sig(772);
CN_in_sig(1801)	<=	VN_out_sig(773);
CN_in_sig(3273)	<=	VN_out_sig(774);
CN_in_sig(4865)	<=	VN_out_sig(775);
CN_in_sig(1089)	<=	VN_out_sig(776);
CN_in_sig(1809)	<=	VN_out_sig(777);
CN_in_sig(3281)	<=	VN_out_sig(778);
CN_in_sig(4873)	<=	VN_out_sig(779);
CN_in_sig(1097)	<=	VN_out_sig(780);
CN_in_sig(1817)	<=	VN_out_sig(781);
CN_in_sig(3289)	<=	VN_out_sig(782);
CN_in_sig(4881)	<=	VN_out_sig(783);
CN_in_sig(1105)	<=	VN_out_sig(784);
CN_in_sig(1825)	<=	VN_out_sig(785);
CN_in_sig(3297)	<=	VN_out_sig(786);
CN_in_sig(4889)	<=	VN_out_sig(787);
CN_in_sig(1113)	<=	VN_out_sig(788);
CN_in_sig(1833)	<=	VN_out_sig(789);
CN_in_sig(3305)	<=	VN_out_sig(790);
CN_in_sig(4897)	<=	VN_out_sig(791);
CN_in_sig(1121)	<=	VN_out_sig(792);
CN_in_sig(1841)	<=	VN_out_sig(793);
CN_in_sig(3313)	<=	VN_out_sig(794);
CN_in_sig(4905)	<=	VN_out_sig(795);
CN_in_sig(1129)	<=	VN_out_sig(796);
CN_in_sig(1849)	<=	VN_out_sig(797);
CN_in_sig(3321)	<=	VN_out_sig(798);
CN_in_sig(4913)	<=	VN_out_sig(799);
CN_in_sig(1137)	<=	VN_out_sig(800);
CN_in_sig(1857)	<=	VN_out_sig(801);
CN_in_sig(3329)	<=	VN_out_sig(802);
CN_in_sig(4921)	<=	VN_out_sig(803);
CN_in_sig(1145)	<=	VN_out_sig(804);
CN_in_sig(1865)	<=	VN_out_sig(805);
CN_in_sig(3337)	<=	VN_out_sig(806);
CN_in_sig(4929)	<=	VN_out_sig(807);
CN_in_sig(1153)	<=	VN_out_sig(808);
CN_in_sig(1873)	<=	VN_out_sig(809);
CN_in_sig(3345)	<=	VN_out_sig(810);
CN_in_sig(4937)	<=	VN_out_sig(811);
CN_in_sig(1161)	<=	VN_out_sig(812);
CN_in_sig(1881)	<=	VN_out_sig(813);
CN_in_sig(3353)	<=	VN_out_sig(814);
CN_in_sig(4945)	<=	VN_out_sig(815);
CN_in_sig(1169)	<=	VN_out_sig(816);
CN_in_sig(1889)	<=	VN_out_sig(817);
CN_in_sig(3361)	<=	VN_out_sig(818);
CN_in_sig(4953)	<=	VN_out_sig(819);
CN_in_sig(1177)	<=	VN_out_sig(820);
CN_in_sig(1897)	<=	VN_out_sig(821);
CN_in_sig(3369)	<=	VN_out_sig(822);
CN_in_sig(4961)	<=	VN_out_sig(823);
CN_in_sig(1185)	<=	VN_out_sig(824);
CN_in_sig(1905)	<=	VN_out_sig(825);
CN_in_sig(3377)	<=	VN_out_sig(826);
CN_in_sig(4969)	<=	VN_out_sig(827);
CN_in_sig(1193)	<=	VN_out_sig(828);
CN_in_sig(1913)	<=	VN_out_sig(829);
CN_in_sig(3385)	<=	VN_out_sig(830);
CN_in_sig(4977)	<=	VN_out_sig(831);
CN_in_sig(1201)	<=	VN_out_sig(832);
CN_in_sig(1921)	<=	VN_out_sig(833);
CN_in_sig(3393)	<=	VN_out_sig(834);
CN_in_sig(4985)	<=	VN_out_sig(835);
CN_in_sig(1209)	<=	VN_out_sig(836);
CN_in_sig(1929)	<=	VN_out_sig(837);
CN_in_sig(3401)	<=	VN_out_sig(838);
CN_in_sig(4993)	<=	VN_out_sig(839);
CN_in_sig(1217)	<=	VN_out_sig(840);
CN_in_sig(1937)	<=	VN_out_sig(841);
CN_in_sig(3409)	<=	VN_out_sig(842);
CN_in_sig(5001)	<=	VN_out_sig(843);
CN_in_sig(1225)	<=	VN_out_sig(844);
CN_in_sig(1945)	<=	VN_out_sig(845);
CN_in_sig(3417)	<=	VN_out_sig(846);
CN_in_sig(5009)	<=	VN_out_sig(847);
CN_in_sig(1233)	<=	VN_out_sig(848);
CN_in_sig(1953)	<=	VN_out_sig(849);
CN_in_sig(3425)	<=	VN_out_sig(850);
CN_in_sig(5017)	<=	VN_out_sig(851);
CN_in_sig(1241)	<=	VN_out_sig(852);
CN_in_sig(1961)	<=	VN_out_sig(853);
CN_in_sig(3433)	<=	VN_out_sig(854);
CN_in_sig(5025)	<=	VN_out_sig(855);
CN_in_sig(1249)	<=	VN_out_sig(856);
CN_in_sig(1969)	<=	VN_out_sig(857);
CN_in_sig(3441)	<=	VN_out_sig(858);
CN_in_sig(5033)	<=	VN_out_sig(859);
CN_in_sig(1257)	<=	VN_out_sig(860);
CN_in_sig(1977)	<=	VN_out_sig(861);
CN_in_sig(3449)	<=	VN_out_sig(862);
CN_in_sig(5041)	<=	VN_out_sig(863);
CN_in_sig(217)	<=	VN_out_sig(864);
CN_in_sig(1457)	<=	VN_out_sig(865);
CN_in_sig(3833)	<=	VN_out_sig(866);
CN_in_sig(4721)	<=	VN_out_sig(867);
CN_in_sig(225)	<=	VN_out_sig(868);
CN_in_sig(1465)	<=	VN_out_sig(869);
CN_in_sig(3841)	<=	VN_out_sig(870);
CN_in_sig(4729)	<=	VN_out_sig(871);
CN_in_sig(233)	<=	VN_out_sig(872);
CN_in_sig(1473)	<=	VN_out_sig(873);
CN_in_sig(3849)	<=	VN_out_sig(874);
CN_in_sig(4737)	<=	VN_out_sig(875);
CN_in_sig(241)	<=	VN_out_sig(876);
CN_in_sig(1481)	<=	VN_out_sig(877);
CN_in_sig(3857)	<=	VN_out_sig(878);
CN_in_sig(4745)	<=	VN_out_sig(879);
CN_in_sig(249)	<=	VN_out_sig(880);
CN_in_sig(1489)	<=	VN_out_sig(881);
CN_in_sig(3865)	<=	VN_out_sig(882);
CN_in_sig(4321)	<=	VN_out_sig(883);
CN_in_sig(257)	<=	VN_out_sig(884);
CN_in_sig(1497)	<=	VN_out_sig(885);
CN_in_sig(3873)	<=	VN_out_sig(886);
CN_in_sig(4329)	<=	VN_out_sig(887);
CN_in_sig(265)	<=	VN_out_sig(888);
CN_in_sig(1505)	<=	VN_out_sig(889);
CN_in_sig(3881)	<=	VN_out_sig(890);
CN_in_sig(4337)	<=	VN_out_sig(891);
CN_in_sig(273)	<=	VN_out_sig(892);
CN_in_sig(1513)	<=	VN_out_sig(893);
CN_in_sig(3457)	<=	VN_out_sig(894);
CN_in_sig(4345)	<=	VN_out_sig(895);
CN_in_sig(281)	<=	VN_out_sig(896);
CN_in_sig(1521)	<=	VN_out_sig(897);
CN_in_sig(3465)	<=	VN_out_sig(898);
CN_in_sig(4353)	<=	VN_out_sig(899);
CN_in_sig(289)	<=	VN_out_sig(900);
CN_in_sig(1529)	<=	VN_out_sig(901);
CN_in_sig(3473)	<=	VN_out_sig(902);
CN_in_sig(4361)	<=	VN_out_sig(903);
CN_in_sig(297)	<=	VN_out_sig(904);
CN_in_sig(1537)	<=	VN_out_sig(905);
CN_in_sig(3481)	<=	VN_out_sig(906);
CN_in_sig(4369)	<=	VN_out_sig(907);
CN_in_sig(305)	<=	VN_out_sig(908);
CN_in_sig(1545)	<=	VN_out_sig(909);
CN_in_sig(3489)	<=	VN_out_sig(910);
CN_in_sig(4377)	<=	VN_out_sig(911);
CN_in_sig(313)	<=	VN_out_sig(912);
CN_in_sig(1553)	<=	VN_out_sig(913);
CN_in_sig(3497)	<=	VN_out_sig(914);
CN_in_sig(4385)	<=	VN_out_sig(915);
CN_in_sig(321)	<=	VN_out_sig(916);
CN_in_sig(1561)	<=	VN_out_sig(917);
CN_in_sig(3505)	<=	VN_out_sig(918);
CN_in_sig(4393)	<=	VN_out_sig(919);
CN_in_sig(329)	<=	VN_out_sig(920);
CN_in_sig(1569)	<=	VN_out_sig(921);
CN_in_sig(3513)	<=	VN_out_sig(922);
CN_in_sig(4401)	<=	VN_out_sig(923);
CN_in_sig(337)	<=	VN_out_sig(924);
CN_in_sig(1577)	<=	VN_out_sig(925);
CN_in_sig(3521)	<=	VN_out_sig(926);
CN_in_sig(4409)	<=	VN_out_sig(927);
CN_in_sig(345)	<=	VN_out_sig(928);
CN_in_sig(1585)	<=	VN_out_sig(929);
CN_in_sig(3529)	<=	VN_out_sig(930);
CN_in_sig(4417)	<=	VN_out_sig(931);
CN_in_sig(353)	<=	VN_out_sig(932);
CN_in_sig(1593)	<=	VN_out_sig(933);
CN_in_sig(3537)	<=	VN_out_sig(934);
CN_in_sig(4425)	<=	VN_out_sig(935);
CN_in_sig(361)	<=	VN_out_sig(936);
CN_in_sig(1601)	<=	VN_out_sig(937);
CN_in_sig(3545)	<=	VN_out_sig(938);
CN_in_sig(4433)	<=	VN_out_sig(939);
CN_in_sig(369)	<=	VN_out_sig(940);
CN_in_sig(1609)	<=	VN_out_sig(941);
CN_in_sig(3553)	<=	VN_out_sig(942);
CN_in_sig(4441)	<=	VN_out_sig(943);
CN_in_sig(377)	<=	VN_out_sig(944);
CN_in_sig(1617)	<=	VN_out_sig(945);
CN_in_sig(3561)	<=	VN_out_sig(946);
CN_in_sig(4449)	<=	VN_out_sig(947);
CN_in_sig(385)	<=	VN_out_sig(948);
CN_in_sig(1625)	<=	VN_out_sig(949);
CN_in_sig(3569)	<=	VN_out_sig(950);
CN_in_sig(4457)	<=	VN_out_sig(951);
CN_in_sig(393)	<=	VN_out_sig(952);
CN_in_sig(1633)	<=	VN_out_sig(953);
CN_in_sig(3577)	<=	VN_out_sig(954);
CN_in_sig(4465)	<=	VN_out_sig(955);
CN_in_sig(401)	<=	VN_out_sig(956);
CN_in_sig(1641)	<=	VN_out_sig(957);
CN_in_sig(3585)	<=	VN_out_sig(958);
CN_in_sig(4473)	<=	VN_out_sig(959);
CN_in_sig(409)	<=	VN_out_sig(960);
CN_in_sig(1649)	<=	VN_out_sig(961);
CN_in_sig(3593)	<=	VN_out_sig(962);
CN_in_sig(4481)	<=	VN_out_sig(963);
CN_in_sig(417)	<=	VN_out_sig(964);
CN_in_sig(1657)	<=	VN_out_sig(965);
CN_in_sig(3601)	<=	VN_out_sig(966);
CN_in_sig(4489)	<=	VN_out_sig(967);
CN_in_sig(425)	<=	VN_out_sig(968);
CN_in_sig(1665)	<=	VN_out_sig(969);
CN_in_sig(3609)	<=	VN_out_sig(970);
CN_in_sig(4497)	<=	VN_out_sig(971);
CN_in_sig(1)	<=	VN_out_sig(972);
CN_in_sig(1673)	<=	VN_out_sig(973);
CN_in_sig(3617)	<=	VN_out_sig(974);
CN_in_sig(4505)	<=	VN_out_sig(975);
CN_in_sig(9)	<=	VN_out_sig(976);
CN_in_sig(1681)	<=	VN_out_sig(977);
CN_in_sig(3625)	<=	VN_out_sig(978);
CN_in_sig(4513)	<=	VN_out_sig(979);
CN_in_sig(17)	<=	VN_out_sig(980);
CN_in_sig(1689)	<=	VN_out_sig(981);
CN_in_sig(3633)	<=	VN_out_sig(982);
CN_in_sig(4521)	<=	VN_out_sig(983);
CN_in_sig(25)	<=	VN_out_sig(984);
CN_in_sig(1697)	<=	VN_out_sig(985);
CN_in_sig(3641)	<=	VN_out_sig(986);
CN_in_sig(4529)	<=	VN_out_sig(987);
CN_in_sig(33)	<=	VN_out_sig(988);
CN_in_sig(1705)	<=	VN_out_sig(989);
CN_in_sig(3649)	<=	VN_out_sig(990);
CN_in_sig(4537)	<=	VN_out_sig(991);
CN_in_sig(41)	<=	VN_out_sig(992);
CN_in_sig(1713)	<=	VN_out_sig(993);
CN_in_sig(3657)	<=	VN_out_sig(994);
CN_in_sig(4545)	<=	VN_out_sig(995);
CN_in_sig(49)	<=	VN_out_sig(996);
CN_in_sig(1721)	<=	VN_out_sig(997);
CN_in_sig(3665)	<=	VN_out_sig(998);
CN_in_sig(4553)	<=	VN_out_sig(999);
CN_in_sig(57)	<=	VN_out_sig(1000);
CN_in_sig(1297)	<=	VN_out_sig(1001);
CN_in_sig(3673)	<=	VN_out_sig(1002);
CN_in_sig(4561)	<=	VN_out_sig(1003);
CN_in_sig(65)	<=	VN_out_sig(1004);
CN_in_sig(1305)	<=	VN_out_sig(1005);
CN_in_sig(3681)	<=	VN_out_sig(1006);
CN_in_sig(4569)	<=	VN_out_sig(1007);
CN_in_sig(73)	<=	VN_out_sig(1008);
CN_in_sig(1313)	<=	VN_out_sig(1009);
CN_in_sig(3689)	<=	VN_out_sig(1010);
CN_in_sig(4577)	<=	VN_out_sig(1011);
CN_in_sig(81)	<=	VN_out_sig(1012);
CN_in_sig(1321)	<=	VN_out_sig(1013);
CN_in_sig(3697)	<=	VN_out_sig(1014);
CN_in_sig(4585)	<=	VN_out_sig(1015);
CN_in_sig(89)	<=	VN_out_sig(1016);
CN_in_sig(1329)	<=	VN_out_sig(1017);
CN_in_sig(3705)	<=	VN_out_sig(1018);
CN_in_sig(4593)	<=	VN_out_sig(1019);
CN_in_sig(97)	<=	VN_out_sig(1020);
CN_in_sig(1337)	<=	VN_out_sig(1021);
CN_in_sig(3713)	<=	VN_out_sig(1022);
CN_in_sig(4601)	<=	VN_out_sig(1023);
CN_in_sig(105)	<=	VN_out_sig(1024);
CN_in_sig(1345)	<=	VN_out_sig(1025);
CN_in_sig(3721)	<=	VN_out_sig(1026);
CN_in_sig(4609)	<=	VN_out_sig(1027);
CN_in_sig(113)	<=	VN_out_sig(1028);
CN_in_sig(1353)	<=	VN_out_sig(1029);
CN_in_sig(3729)	<=	VN_out_sig(1030);
CN_in_sig(4617)	<=	VN_out_sig(1031);
CN_in_sig(121)	<=	VN_out_sig(1032);
CN_in_sig(1361)	<=	VN_out_sig(1033);
CN_in_sig(3737)	<=	VN_out_sig(1034);
CN_in_sig(4625)	<=	VN_out_sig(1035);
CN_in_sig(129)	<=	VN_out_sig(1036);
CN_in_sig(1369)	<=	VN_out_sig(1037);
CN_in_sig(3745)	<=	VN_out_sig(1038);
CN_in_sig(4633)	<=	VN_out_sig(1039);
CN_in_sig(137)	<=	VN_out_sig(1040);
CN_in_sig(1377)	<=	VN_out_sig(1041);
CN_in_sig(3753)	<=	VN_out_sig(1042);
CN_in_sig(4641)	<=	VN_out_sig(1043);
CN_in_sig(145)	<=	VN_out_sig(1044);
CN_in_sig(1385)	<=	VN_out_sig(1045);
CN_in_sig(3761)	<=	VN_out_sig(1046);
CN_in_sig(4649)	<=	VN_out_sig(1047);
CN_in_sig(153)	<=	VN_out_sig(1048);
CN_in_sig(1393)	<=	VN_out_sig(1049);
CN_in_sig(3769)	<=	VN_out_sig(1050);
CN_in_sig(4657)	<=	VN_out_sig(1051);
CN_in_sig(161)	<=	VN_out_sig(1052);
CN_in_sig(1401)	<=	VN_out_sig(1053);
CN_in_sig(3777)	<=	VN_out_sig(1054);
CN_in_sig(4665)	<=	VN_out_sig(1055);
CN_in_sig(169)	<=	VN_out_sig(1056);
CN_in_sig(1409)	<=	VN_out_sig(1057);
CN_in_sig(3785)	<=	VN_out_sig(1058);
CN_in_sig(4673)	<=	VN_out_sig(1059);
CN_in_sig(177)	<=	VN_out_sig(1060);
CN_in_sig(1417)	<=	VN_out_sig(1061);
CN_in_sig(3793)	<=	VN_out_sig(1062);
CN_in_sig(4681)	<=	VN_out_sig(1063);
CN_in_sig(185)	<=	VN_out_sig(1064);
CN_in_sig(1425)	<=	VN_out_sig(1065);
CN_in_sig(3801)	<=	VN_out_sig(1066);
CN_in_sig(4689)	<=	VN_out_sig(1067);
CN_in_sig(193)	<=	VN_out_sig(1068);
CN_in_sig(1433)	<=	VN_out_sig(1069);
CN_in_sig(3809)	<=	VN_out_sig(1070);
CN_in_sig(4697)	<=	VN_out_sig(1071);
CN_in_sig(201)	<=	VN_out_sig(1072);
CN_in_sig(1441)	<=	VN_out_sig(1073);
CN_in_sig(3817)	<=	VN_out_sig(1074);
CN_in_sig(4705)	<=	VN_out_sig(1075);
CN_in_sig(209)	<=	VN_out_sig(1076);
CN_in_sig(1449)	<=	VN_out_sig(1077);
CN_in_sig(3825)	<=	VN_out_sig(1078);
CN_in_sig(4713)	<=	VN_out_sig(1079);
CN_in_sig(617)	<=	VN_out_sig(1080);
CN_in_sig(2513)	<=	VN_out_sig(1081);
CN_in_sig(2745)	<=	VN_out_sig(1082);
CN_in_sig(4297)	<=	VN_out_sig(1083);
CN_in_sig(625)	<=	VN_out_sig(1084);
CN_in_sig(2521)	<=	VN_out_sig(1085);
CN_in_sig(2753)	<=	VN_out_sig(1086);
CN_in_sig(4305)	<=	VN_out_sig(1087);
CN_in_sig(633)	<=	VN_out_sig(1088);
CN_in_sig(2529)	<=	VN_out_sig(1089);
CN_in_sig(2761)	<=	VN_out_sig(1090);
CN_in_sig(4313)	<=	VN_out_sig(1091);
CN_in_sig(641)	<=	VN_out_sig(1092);
CN_in_sig(2537)	<=	VN_out_sig(1093);
CN_in_sig(2769)	<=	VN_out_sig(1094);
CN_in_sig(3889)	<=	VN_out_sig(1095);
CN_in_sig(649)	<=	VN_out_sig(1096);
CN_in_sig(2545)	<=	VN_out_sig(1097);
CN_in_sig(2777)	<=	VN_out_sig(1098);
CN_in_sig(3897)	<=	VN_out_sig(1099);
CN_in_sig(657)	<=	VN_out_sig(1100);
CN_in_sig(2553)	<=	VN_out_sig(1101);
CN_in_sig(2785)	<=	VN_out_sig(1102);
CN_in_sig(3905)	<=	VN_out_sig(1103);
CN_in_sig(665)	<=	VN_out_sig(1104);
CN_in_sig(2561)	<=	VN_out_sig(1105);
CN_in_sig(2793)	<=	VN_out_sig(1106);
CN_in_sig(3913)	<=	VN_out_sig(1107);
CN_in_sig(673)	<=	VN_out_sig(1108);
CN_in_sig(2569)	<=	VN_out_sig(1109);
CN_in_sig(2801)	<=	VN_out_sig(1110);
CN_in_sig(3921)	<=	VN_out_sig(1111);
CN_in_sig(681)	<=	VN_out_sig(1112);
CN_in_sig(2577)	<=	VN_out_sig(1113);
CN_in_sig(2809)	<=	VN_out_sig(1114);
CN_in_sig(3929)	<=	VN_out_sig(1115);
CN_in_sig(689)	<=	VN_out_sig(1116);
CN_in_sig(2585)	<=	VN_out_sig(1117);
CN_in_sig(2817)	<=	VN_out_sig(1118);
CN_in_sig(3937)	<=	VN_out_sig(1119);
CN_in_sig(697)	<=	VN_out_sig(1120);
CN_in_sig(2161)	<=	VN_out_sig(1121);
CN_in_sig(2825)	<=	VN_out_sig(1122);
CN_in_sig(3945)	<=	VN_out_sig(1123);
CN_in_sig(705)	<=	VN_out_sig(1124);
CN_in_sig(2169)	<=	VN_out_sig(1125);
CN_in_sig(2833)	<=	VN_out_sig(1126);
CN_in_sig(3953)	<=	VN_out_sig(1127);
CN_in_sig(713)	<=	VN_out_sig(1128);
CN_in_sig(2177)	<=	VN_out_sig(1129);
CN_in_sig(2841)	<=	VN_out_sig(1130);
CN_in_sig(3961)	<=	VN_out_sig(1131);
CN_in_sig(721)	<=	VN_out_sig(1132);
CN_in_sig(2185)	<=	VN_out_sig(1133);
CN_in_sig(2849)	<=	VN_out_sig(1134);
CN_in_sig(3969)	<=	VN_out_sig(1135);
CN_in_sig(729)	<=	VN_out_sig(1136);
CN_in_sig(2193)	<=	VN_out_sig(1137);
CN_in_sig(2857)	<=	VN_out_sig(1138);
CN_in_sig(3977)	<=	VN_out_sig(1139);
CN_in_sig(737)	<=	VN_out_sig(1140);
CN_in_sig(2201)	<=	VN_out_sig(1141);
CN_in_sig(2865)	<=	VN_out_sig(1142);
CN_in_sig(3985)	<=	VN_out_sig(1143);
CN_in_sig(745)	<=	VN_out_sig(1144);
CN_in_sig(2209)	<=	VN_out_sig(1145);
CN_in_sig(2873)	<=	VN_out_sig(1146);
CN_in_sig(3993)	<=	VN_out_sig(1147);
CN_in_sig(753)	<=	VN_out_sig(1148);
CN_in_sig(2217)	<=	VN_out_sig(1149);
CN_in_sig(2881)	<=	VN_out_sig(1150);
CN_in_sig(4001)	<=	VN_out_sig(1151);
CN_in_sig(761)	<=	VN_out_sig(1152);
CN_in_sig(2225)	<=	VN_out_sig(1153);
CN_in_sig(2889)	<=	VN_out_sig(1154);
CN_in_sig(4009)	<=	VN_out_sig(1155);
CN_in_sig(769)	<=	VN_out_sig(1156);
CN_in_sig(2233)	<=	VN_out_sig(1157);
CN_in_sig(2897)	<=	VN_out_sig(1158);
CN_in_sig(4017)	<=	VN_out_sig(1159);
CN_in_sig(777)	<=	VN_out_sig(1160);
CN_in_sig(2241)	<=	VN_out_sig(1161);
CN_in_sig(2905)	<=	VN_out_sig(1162);
CN_in_sig(4025)	<=	VN_out_sig(1163);
CN_in_sig(785)	<=	VN_out_sig(1164);
CN_in_sig(2249)	<=	VN_out_sig(1165);
CN_in_sig(2913)	<=	VN_out_sig(1166);
CN_in_sig(4033)	<=	VN_out_sig(1167);
CN_in_sig(793)	<=	VN_out_sig(1168);
CN_in_sig(2257)	<=	VN_out_sig(1169);
CN_in_sig(2921)	<=	VN_out_sig(1170);
CN_in_sig(4041)	<=	VN_out_sig(1171);
CN_in_sig(801)	<=	VN_out_sig(1172);
CN_in_sig(2265)	<=	VN_out_sig(1173);
CN_in_sig(2929)	<=	VN_out_sig(1174);
CN_in_sig(4049)	<=	VN_out_sig(1175);
CN_in_sig(809)	<=	VN_out_sig(1176);
CN_in_sig(2273)	<=	VN_out_sig(1177);
CN_in_sig(2937)	<=	VN_out_sig(1178);
CN_in_sig(4057)	<=	VN_out_sig(1179);
CN_in_sig(817)	<=	VN_out_sig(1180);
CN_in_sig(2281)	<=	VN_out_sig(1181);
CN_in_sig(2945)	<=	VN_out_sig(1182);
CN_in_sig(4065)	<=	VN_out_sig(1183);
CN_in_sig(825)	<=	VN_out_sig(1184);
CN_in_sig(2289)	<=	VN_out_sig(1185);
CN_in_sig(2953)	<=	VN_out_sig(1186);
CN_in_sig(4073)	<=	VN_out_sig(1187);
CN_in_sig(833)	<=	VN_out_sig(1188);
CN_in_sig(2297)	<=	VN_out_sig(1189);
CN_in_sig(2961)	<=	VN_out_sig(1190);
CN_in_sig(4081)	<=	VN_out_sig(1191);
CN_in_sig(841)	<=	VN_out_sig(1192);
CN_in_sig(2305)	<=	VN_out_sig(1193);
CN_in_sig(2969)	<=	VN_out_sig(1194);
CN_in_sig(4089)	<=	VN_out_sig(1195);
CN_in_sig(849)	<=	VN_out_sig(1196);
CN_in_sig(2313)	<=	VN_out_sig(1197);
CN_in_sig(2977)	<=	VN_out_sig(1198);
CN_in_sig(4097)	<=	VN_out_sig(1199);
CN_in_sig(857)	<=	VN_out_sig(1200);
CN_in_sig(2321)	<=	VN_out_sig(1201);
CN_in_sig(2985)	<=	VN_out_sig(1202);
CN_in_sig(4105)	<=	VN_out_sig(1203);
CN_in_sig(433)	<=	VN_out_sig(1204);
CN_in_sig(2329)	<=	VN_out_sig(1205);
CN_in_sig(2993)	<=	VN_out_sig(1206);
CN_in_sig(4113)	<=	VN_out_sig(1207);
CN_in_sig(441)	<=	VN_out_sig(1208);
CN_in_sig(2337)	<=	VN_out_sig(1209);
CN_in_sig(3001)	<=	VN_out_sig(1210);
CN_in_sig(4121)	<=	VN_out_sig(1211);
CN_in_sig(449)	<=	VN_out_sig(1212);
CN_in_sig(2345)	<=	VN_out_sig(1213);
CN_in_sig(3009)	<=	VN_out_sig(1214);
CN_in_sig(4129)	<=	VN_out_sig(1215);
CN_in_sig(457)	<=	VN_out_sig(1216);
CN_in_sig(2353)	<=	VN_out_sig(1217);
CN_in_sig(3017)	<=	VN_out_sig(1218);
CN_in_sig(4137)	<=	VN_out_sig(1219);
CN_in_sig(465)	<=	VN_out_sig(1220);
CN_in_sig(2361)	<=	VN_out_sig(1221);
CN_in_sig(2593)	<=	VN_out_sig(1222);
CN_in_sig(4145)	<=	VN_out_sig(1223);
CN_in_sig(473)	<=	VN_out_sig(1224);
CN_in_sig(2369)	<=	VN_out_sig(1225);
CN_in_sig(2601)	<=	VN_out_sig(1226);
CN_in_sig(4153)	<=	VN_out_sig(1227);
CN_in_sig(481)	<=	VN_out_sig(1228);
CN_in_sig(2377)	<=	VN_out_sig(1229);
CN_in_sig(2609)	<=	VN_out_sig(1230);
CN_in_sig(4161)	<=	VN_out_sig(1231);
CN_in_sig(489)	<=	VN_out_sig(1232);
CN_in_sig(2385)	<=	VN_out_sig(1233);
CN_in_sig(2617)	<=	VN_out_sig(1234);
CN_in_sig(4169)	<=	VN_out_sig(1235);
CN_in_sig(497)	<=	VN_out_sig(1236);
CN_in_sig(2393)	<=	VN_out_sig(1237);
CN_in_sig(2625)	<=	VN_out_sig(1238);
CN_in_sig(4177)	<=	VN_out_sig(1239);
CN_in_sig(505)	<=	VN_out_sig(1240);
CN_in_sig(2401)	<=	VN_out_sig(1241);
CN_in_sig(2633)	<=	VN_out_sig(1242);
CN_in_sig(4185)	<=	VN_out_sig(1243);
CN_in_sig(513)	<=	VN_out_sig(1244);
CN_in_sig(2409)	<=	VN_out_sig(1245);
CN_in_sig(2641)	<=	VN_out_sig(1246);
CN_in_sig(4193)	<=	VN_out_sig(1247);
CN_in_sig(521)	<=	VN_out_sig(1248);
CN_in_sig(2417)	<=	VN_out_sig(1249);
CN_in_sig(2649)	<=	VN_out_sig(1250);
CN_in_sig(4201)	<=	VN_out_sig(1251);
CN_in_sig(529)	<=	VN_out_sig(1252);
CN_in_sig(2425)	<=	VN_out_sig(1253);
CN_in_sig(2657)	<=	VN_out_sig(1254);
CN_in_sig(4209)	<=	VN_out_sig(1255);
CN_in_sig(537)	<=	VN_out_sig(1256);
CN_in_sig(2433)	<=	VN_out_sig(1257);
CN_in_sig(2665)	<=	VN_out_sig(1258);
CN_in_sig(4217)	<=	VN_out_sig(1259);
CN_in_sig(545)	<=	VN_out_sig(1260);
CN_in_sig(2441)	<=	VN_out_sig(1261);
CN_in_sig(2673)	<=	VN_out_sig(1262);
CN_in_sig(4225)	<=	VN_out_sig(1263);
CN_in_sig(553)	<=	VN_out_sig(1264);
CN_in_sig(2449)	<=	VN_out_sig(1265);
CN_in_sig(2681)	<=	VN_out_sig(1266);
CN_in_sig(4233)	<=	VN_out_sig(1267);
CN_in_sig(561)	<=	VN_out_sig(1268);
CN_in_sig(2457)	<=	VN_out_sig(1269);
CN_in_sig(2689)	<=	VN_out_sig(1270);
CN_in_sig(4241)	<=	VN_out_sig(1271);
CN_in_sig(569)	<=	VN_out_sig(1272);
CN_in_sig(2465)	<=	VN_out_sig(1273);
CN_in_sig(2697)	<=	VN_out_sig(1274);
CN_in_sig(4249)	<=	VN_out_sig(1275);
CN_in_sig(577)	<=	VN_out_sig(1276);
CN_in_sig(2473)	<=	VN_out_sig(1277);
CN_in_sig(2705)	<=	VN_out_sig(1278);
CN_in_sig(4257)	<=	VN_out_sig(1279);
CN_in_sig(585)	<=	VN_out_sig(1280);
CN_in_sig(2481)	<=	VN_out_sig(1281);
CN_in_sig(2713)	<=	VN_out_sig(1282);
CN_in_sig(4265)	<=	VN_out_sig(1283);
CN_in_sig(593)	<=	VN_out_sig(1284);
CN_in_sig(2489)	<=	VN_out_sig(1285);
CN_in_sig(2721)	<=	VN_out_sig(1286);
CN_in_sig(4273)	<=	VN_out_sig(1287);
CN_in_sig(601)	<=	VN_out_sig(1288);
CN_in_sig(2497)	<=	VN_out_sig(1289);
CN_in_sig(2729)	<=	VN_out_sig(1290);
CN_in_sig(4281)	<=	VN_out_sig(1291);
CN_in_sig(609)	<=	VN_out_sig(1292);
CN_in_sig(2505)	<=	VN_out_sig(1293);
CN_in_sig(2737)	<=	VN_out_sig(1294);
CN_in_sig(4289)	<=	VN_out_sig(1295);
CN_in_sig(634)	<=	VN_out_sig(1296);
CN_in_sig(1570)	<=	VN_out_sig(1297);
CN_in_sig(3730)	<=	VN_out_sig(1298);
CN_in_sig(4898)	<=	VN_out_sig(1299);
CN_in_sig(642)	<=	VN_out_sig(1300);
CN_in_sig(1578)	<=	VN_out_sig(1301);
CN_in_sig(3738)	<=	VN_out_sig(1302);
CN_in_sig(4906)	<=	VN_out_sig(1303);
CN_in_sig(650)	<=	VN_out_sig(1304);
CN_in_sig(1586)	<=	VN_out_sig(1305);
CN_in_sig(3746)	<=	VN_out_sig(1306);
CN_in_sig(4914)	<=	VN_out_sig(1307);
CN_in_sig(658)	<=	VN_out_sig(1308);
CN_in_sig(1594)	<=	VN_out_sig(1309);
CN_in_sig(3754)	<=	VN_out_sig(1310);
CN_in_sig(4922)	<=	VN_out_sig(1311);
CN_in_sig(666)	<=	VN_out_sig(1312);
CN_in_sig(1602)	<=	VN_out_sig(1313);
CN_in_sig(3762)	<=	VN_out_sig(1314);
CN_in_sig(4930)	<=	VN_out_sig(1315);
CN_in_sig(674)	<=	VN_out_sig(1316);
CN_in_sig(1610)	<=	VN_out_sig(1317);
CN_in_sig(3770)	<=	VN_out_sig(1318);
CN_in_sig(4938)	<=	VN_out_sig(1319);
CN_in_sig(682)	<=	VN_out_sig(1320);
CN_in_sig(1618)	<=	VN_out_sig(1321);
CN_in_sig(3778)	<=	VN_out_sig(1322);
CN_in_sig(4946)	<=	VN_out_sig(1323);
CN_in_sig(690)	<=	VN_out_sig(1324);
CN_in_sig(1626)	<=	VN_out_sig(1325);
CN_in_sig(3786)	<=	VN_out_sig(1326);
CN_in_sig(4954)	<=	VN_out_sig(1327);
CN_in_sig(698)	<=	VN_out_sig(1328);
CN_in_sig(1634)	<=	VN_out_sig(1329);
CN_in_sig(3794)	<=	VN_out_sig(1330);
CN_in_sig(4962)	<=	VN_out_sig(1331);
CN_in_sig(706)	<=	VN_out_sig(1332);
CN_in_sig(1642)	<=	VN_out_sig(1333);
CN_in_sig(3802)	<=	VN_out_sig(1334);
CN_in_sig(4970)	<=	VN_out_sig(1335);
CN_in_sig(714)	<=	VN_out_sig(1336);
CN_in_sig(1650)	<=	VN_out_sig(1337);
CN_in_sig(3810)	<=	VN_out_sig(1338);
CN_in_sig(4978)	<=	VN_out_sig(1339);
CN_in_sig(722)	<=	VN_out_sig(1340);
CN_in_sig(1658)	<=	VN_out_sig(1341);
CN_in_sig(3818)	<=	VN_out_sig(1342);
CN_in_sig(4986)	<=	VN_out_sig(1343);
CN_in_sig(730)	<=	VN_out_sig(1344);
CN_in_sig(1666)	<=	VN_out_sig(1345);
CN_in_sig(3826)	<=	VN_out_sig(1346);
CN_in_sig(4994)	<=	VN_out_sig(1347);
CN_in_sig(738)	<=	VN_out_sig(1348);
CN_in_sig(1674)	<=	VN_out_sig(1349);
CN_in_sig(3834)	<=	VN_out_sig(1350);
CN_in_sig(5002)	<=	VN_out_sig(1351);
CN_in_sig(746)	<=	VN_out_sig(1352);
CN_in_sig(1682)	<=	VN_out_sig(1353);
CN_in_sig(3842)	<=	VN_out_sig(1354);
CN_in_sig(5010)	<=	VN_out_sig(1355);
CN_in_sig(754)	<=	VN_out_sig(1356);
CN_in_sig(1690)	<=	VN_out_sig(1357);
CN_in_sig(3850)	<=	VN_out_sig(1358);
CN_in_sig(5018)	<=	VN_out_sig(1359);
CN_in_sig(762)	<=	VN_out_sig(1360);
CN_in_sig(1698)	<=	VN_out_sig(1361);
CN_in_sig(3858)	<=	VN_out_sig(1362);
CN_in_sig(5026)	<=	VN_out_sig(1363);
CN_in_sig(770)	<=	VN_out_sig(1364);
CN_in_sig(1706)	<=	VN_out_sig(1365);
CN_in_sig(3866)	<=	VN_out_sig(1366);
CN_in_sig(5034)	<=	VN_out_sig(1367);
CN_in_sig(778)	<=	VN_out_sig(1368);
CN_in_sig(1714)	<=	VN_out_sig(1369);
CN_in_sig(3874)	<=	VN_out_sig(1370);
CN_in_sig(5042)	<=	VN_out_sig(1371);
CN_in_sig(786)	<=	VN_out_sig(1372);
CN_in_sig(1722)	<=	VN_out_sig(1373);
CN_in_sig(3882)	<=	VN_out_sig(1374);
CN_in_sig(5050)	<=	VN_out_sig(1375);
CN_in_sig(794)	<=	VN_out_sig(1376);
CN_in_sig(1298)	<=	VN_out_sig(1377);
CN_in_sig(3458)	<=	VN_out_sig(1378);
CN_in_sig(5058)	<=	VN_out_sig(1379);
CN_in_sig(802)	<=	VN_out_sig(1380);
CN_in_sig(1306)	<=	VN_out_sig(1381);
CN_in_sig(3466)	<=	VN_out_sig(1382);
CN_in_sig(5066)	<=	VN_out_sig(1383);
CN_in_sig(810)	<=	VN_out_sig(1384);
CN_in_sig(1314)	<=	VN_out_sig(1385);
CN_in_sig(3474)	<=	VN_out_sig(1386);
CN_in_sig(5074)	<=	VN_out_sig(1387);
CN_in_sig(818)	<=	VN_out_sig(1388);
CN_in_sig(1322)	<=	VN_out_sig(1389);
CN_in_sig(3482)	<=	VN_out_sig(1390);
CN_in_sig(5082)	<=	VN_out_sig(1391);
CN_in_sig(826)	<=	VN_out_sig(1392);
CN_in_sig(1330)	<=	VN_out_sig(1393);
CN_in_sig(3490)	<=	VN_out_sig(1394);
CN_in_sig(5090)	<=	VN_out_sig(1395);
CN_in_sig(834)	<=	VN_out_sig(1396);
CN_in_sig(1338)	<=	VN_out_sig(1397);
CN_in_sig(3498)	<=	VN_out_sig(1398);
CN_in_sig(5098)	<=	VN_out_sig(1399);
CN_in_sig(842)	<=	VN_out_sig(1400);
CN_in_sig(1346)	<=	VN_out_sig(1401);
CN_in_sig(3506)	<=	VN_out_sig(1402);
CN_in_sig(5106)	<=	VN_out_sig(1403);
CN_in_sig(850)	<=	VN_out_sig(1404);
CN_in_sig(1354)	<=	VN_out_sig(1405);
CN_in_sig(3514)	<=	VN_out_sig(1406);
CN_in_sig(5114)	<=	VN_out_sig(1407);
CN_in_sig(858)	<=	VN_out_sig(1408);
CN_in_sig(1362)	<=	VN_out_sig(1409);
CN_in_sig(3522)	<=	VN_out_sig(1410);
CN_in_sig(5122)	<=	VN_out_sig(1411);
CN_in_sig(434)	<=	VN_out_sig(1412);
CN_in_sig(1370)	<=	VN_out_sig(1413);
CN_in_sig(3530)	<=	VN_out_sig(1414);
CN_in_sig(5130)	<=	VN_out_sig(1415);
CN_in_sig(442)	<=	VN_out_sig(1416);
CN_in_sig(1378)	<=	VN_out_sig(1417);
CN_in_sig(3538)	<=	VN_out_sig(1418);
CN_in_sig(5138)	<=	VN_out_sig(1419);
CN_in_sig(450)	<=	VN_out_sig(1420);
CN_in_sig(1386)	<=	VN_out_sig(1421);
CN_in_sig(3546)	<=	VN_out_sig(1422);
CN_in_sig(5146)	<=	VN_out_sig(1423);
CN_in_sig(458)	<=	VN_out_sig(1424);
CN_in_sig(1394)	<=	VN_out_sig(1425);
CN_in_sig(3554)	<=	VN_out_sig(1426);
CN_in_sig(5154)	<=	VN_out_sig(1427);
CN_in_sig(466)	<=	VN_out_sig(1428);
CN_in_sig(1402)	<=	VN_out_sig(1429);
CN_in_sig(3562)	<=	VN_out_sig(1430);
CN_in_sig(5162)	<=	VN_out_sig(1431);
CN_in_sig(474)	<=	VN_out_sig(1432);
CN_in_sig(1410)	<=	VN_out_sig(1433);
CN_in_sig(3570)	<=	VN_out_sig(1434);
CN_in_sig(5170)	<=	VN_out_sig(1435);
CN_in_sig(482)	<=	VN_out_sig(1436);
CN_in_sig(1418)	<=	VN_out_sig(1437);
CN_in_sig(3578)	<=	VN_out_sig(1438);
CN_in_sig(5178)	<=	VN_out_sig(1439);
CN_in_sig(490)	<=	VN_out_sig(1440);
CN_in_sig(1426)	<=	VN_out_sig(1441);
CN_in_sig(3586)	<=	VN_out_sig(1442);
CN_in_sig(4754)	<=	VN_out_sig(1443);
CN_in_sig(498)	<=	VN_out_sig(1444);
CN_in_sig(1434)	<=	VN_out_sig(1445);
CN_in_sig(3594)	<=	VN_out_sig(1446);
CN_in_sig(4762)	<=	VN_out_sig(1447);
CN_in_sig(506)	<=	VN_out_sig(1448);
CN_in_sig(1442)	<=	VN_out_sig(1449);
CN_in_sig(3602)	<=	VN_out_sig(1450);
CN_in_sig(4770)	<=	VN_out_sig(1451);
CN_in_sig(514)	<=	VN_out_sig(1452);
CN_in_sig(1450)	<=	VN_out_sig(1453);
CN_in_sig(3610)	<=	VN_out_sig(1454);
CN_in_sig(4778)	<=	VN_out_sig(1455);
CN_in_sig(522)	<=	VN_out_sig(1456);
CN_in_sig(1458)	<=	VN_out_sig(1457);
CN_in_sig(3618)	<=	VN_out_sig(1458);
CN_in_sig(4786)	<=	VN_out_sig(1459);
CN_in_sig(530)	<=	VN_out_sig(1460);
CN_in_sig(1466)	<=	VN_out_sig(1461);
CN_in_sig(3626)	<=	VN_out_sig(1462);
CN_in_sig(4794)	<=	VN_out_sig(1463);
CN_in_sig(538)	<=	VN_out_sig(1464);
CN_in_sig(1474)	<=	VN_out_sig(1465);
CN_in_sig(3634)	<=	VN_out_sig(1466);
CN_in_sig(4802)	<=	VN_out_sig(1467);
CN_in_sig(546)	<=	VN_out_sig(1468);
CN_in_sig(1482)	<=	VN_out_sig(1469);
CN_in_sig(3642)	<=	VN_out_sig(1470);
CN_in_sig(4810)	<=	VN_out_sig(1471);
CN_in_sig(554)	<=	VN_out_sig(1472);
CN_in_sig(1490)	<=	VN_out_sig(1473);
CN_in_sig(3650)	<=	VN_out_sig(1474);
CN_in_sig(4818)	<=	VN_out_sig(1475);
CN_in_sig(562)	<=	VN_out_sig(1476);
CN_in_sig(1498)	<=	VN_out_sig(1477);
CN_in_sig(3658)	<=	VN_out_sig(1478);
CN_in_sig(4826)	<=	VN_out_sig(1479);
CN_in_sig(570)	<=	VN_out_sig(1480);
CN_in_sig(1506)	<=	VN_out_sig(1481);
CN_in_sig(3666)	<=	VN_out_sig(1482);
CN_in_sig(4834)	<=	VN_out_sig(1483);
CN_in_sig(578)	<=	VN_out_sig(1484);
CN_in_sig(1514)	<=	VN_out_sig(1485);
CN_in_sig(3674)	<=	VN_out_sig(1486);
CN_in_sig(4842)	<=	VN_out_sig(1487);
CN_in_sig(586)	<=	VN_out_sig(1488);
CN_in_sig(1522)	<=	VN_out_sig(1489);
CN_in_sig(3682)	<=	VN_out_sig(1490);
CN_in_sig(4850)	<=	VN_out_sig(1491);
CN_in_sig(594)	<=	VN_out_sig(1492);
CN_in_sig(1530)	<=	VN_out_sig(1493);
CN_in_sig(3690)	<=	VN_out_sig(1494);
CN_in_sig(4858)	<=	VN_out_sig(1495);
CN_in_sig(602)	<=	VN_out_sig(1496);
CN_in_sig(1538)	<=	VN_out_sig(1497);
CN_in_sig(3698)	<=	VN_out_sig(1498);
CN_in_sig(4866)	<=	VN_out_sig(1499);
CN_in_sig(610)	<=	VN_out_sig(1500);
CN_in_sig(1546)	<=	VN_out_sig(1501);
CN_in_sig(3706)	<=	VN_out_sig(1502);
CN_in_sig(4874)	<=	VN_out_sig(1503);
CN_in_sig(618)	<=	VN_out_sig(1504);
CN_in_sig(1554)	<=	VN_out_sig(1505);
CN_in_sig(3714)	<=	VN_out_sig(1506);
CN_in_sig(4882)	<=	VN_out_sig(1507);
CN_in_sig(626)	<=	VN_out_sig(1508);
CN_in_sig(1562)	<=	VN_out_sig(1509);
CN_in_sig(3722)	<=	VN_out_sig(1510);
CN_in_sig(4890)	<=	VN_out_sig(1511);
CN_in_sig(1210)	<=	VN_out_sig(1512);
CN_in_sig(2074)	<=	VN_out_sig(1513);
CN_in_sig(3226)	<=	VN_out_sig(1514);
CN_in_sig(4714)	<=	VN_out_sig(1515);
CN_in_sig(1218)	<=	VN_out_sig(1516);
CN_in_sig(2082)	<=	VN_out_sig(1517);
CN_in_sig(3234)	<=	VN_out_sig(1518);
CN_in_sig(4722)	<=	VN_out_sig(1519);
CN_in_sig(1226)	<=	VN_out_sig(1520);
CN_in_sig(2090)	<=	VN_out_sig(1521);
CN_in_sig(3242)	<=	VN_out_sig(1522);
CN_in_sig(4730)	<=	VN_out_sig(1523);
CN_in_sig(1234)	<=	VN_out_sig(1524);
CN_in_sig(2098)	<=	VN_out_sig(1525);
CN_in_sig(3250)	<=	VN_out_sig(1526);
CN_in_sig(4738)	<=	VN_out_sig(1527);
CN_in_sig(1242)	<=	VN_out_sig(1528);
CN_in_sig(2106)	<=	VN_out_sig(1529);
CN_in_sig(3258)	<=	VN_out_sig(1530);
CN_in_sig(4746)	<=	VN_out_sig(1531);
CN_in_sig(1250)	<=	VN_out_sig(1532);
CN_in_sig(2114)	<=	VN_out_sig(1533);
CN_in_sig(3266)	<=	VN_out_sig(1534);
CN_in_sig(4322)	<=	VN_out_sig(1535);
CN_in_sig(1258)	<=	VN_out_sig(1536);
CN_in_sig(2122)	<=	VN_out_sig(1537);
CN_in_sig(3274)	<=	VN_out_sig(1538);
CN_in_sig(4330)	<=	VN_out_sig(1539);
CN_in_sig(1266)	<=	VN_out_sig(1540);
CN_in_sig(2130)	<=	VN_out_sig(1541);
CN_in_sig(3282)	<=	VN_out_sig(1542);
CN_in_sig(4338)	<=	VN_out_sig(1543);
CN_in_sig(1274)	<=	VN_out_sig(1544);
CN_in_sig(2138)	<=	VN_out_sig(1545);
CN_in_sig(3290)	<=	VN_out_sig(1546);
CN_in_sig(4346)	<=	VN_out_sig(1547);
CN_in_sig(1282)	<=	VN_out_sig(1548);
CN_in_sig(2146)	<=	VN_out_sig(1549);
CN_in_sig(3298)	<=	VN_out_sig(1550);
CN_in_sig(4354)	<=	VN_out_sig(1551);
CN_in_sig(1290)	<=	VN_out_sig(1552);
CN_in_sig(2154)	<=	VN_out_sig(1553);
CN_in_sig(3306)	<=	VN_out_sig(1554);
CN_in_sig(4362)	<=	VN_out_sig(1555);
CN_in_sig(866)	<=	VN_out_sig(1556);
CN_in_sig(1730)	<=	VN_out_sig(1557);
CN_in_sig(3314)	<=	VN_out_sig(1558);
CN_in_sig(4370)	<=	VN_out_sig(1559);
CN_in_sig(874)	<=	VN_out_sig(1560);
CN_in_sig(1738)	<=	VN_out_sig(1561);
CN_in_sig(3322)	<=	VN_out_sig(1562);
CN_in_sig(4378)	<=	VN_out_sig(1563);
CN_in_sig(882)	<=	VN_out_sig(1564);
CN_in_sig(1746)	<=	VN_out_sig(1565);
CN_in_sig(3330)	<=	VN_out_sig(1566);
CN_in_sig(4386)	<=	VN_out_sig(1567);
CN_in_sig(890)	<=	VN_out_sig(1568);
CN_in_sig(1754)	<=	VN_out_sig(1569);
CN_in_sig(3338)	<=	VN_out_sig(1570);
CN_in_sig(4394)	<=	VN_out_sig(1571);
CN_in_sig(898)	<=	VN_out_sig(1572);
CN_in_sig(1762)	<=	VN_out_sig(1573);
CN_in_sig(3346)	<=	VN_out_sig(1574);
CN_in_sig(4402)	<=	VN_out_sig(1575);
CN_in_sig(906)	<=	VN_out_sig(1576);
CN_in_sig(1770)	<=	VN_out_sig(1577);
CN_in_sig(3354)	<=	VN_out_sig(1578);
CN_in_sig(4410)	<=	VN_out_sig(1579);
CN_in_sig(914)	<=	VN_out_sig(1580);
CN_in_sig(1778)	<=	VN_out_sig(1581);
CN_in_sig(3362)	<=	VN_out_sig(1582);
CN_in_sig(4418)	<=	VN_out_sig(1583);
CN_in_sig(922)	<=	VN_out_sig(1584);
CN_in_sig(1786)	<=	VN_out_sig(1585);
CN_in_sig(3370)	<=	VN_out_sig(1586);
CN_in_sig(4426)	<=	VN_out_sig(1587);
CN_in_sig(930)	<=	VN_out_sig(1588);
CN_in_sig(1794)	<=	VN_out_sig(1589);
CN_in_sig(3378)	<=	VN_out_sig(1590);
CN_in_sig(4434)	<=	VN_out_sig(1591);
CN_in_sig(938)	<=	VN_out_sig(1592);
CN_in_sig(1802)	<=	VN_out_sig(1593);
CN_in_sig(3386)	<=	VN_out_sig(1594);
CN_in_sig(4442)	<=	VN_out_sig(1595);
CN_in_sig(946)	<=	VN_out_sig(1596);
CN_in_sig(1810)	<=	VN_out_sig(1597);
CN_in_sig(3394)	<=	VN_out_sig(1598);
CN_in_sig(4450)	<=	VN_out_sig(1599);
CN_in_sig(954)	<=	VN_out_sig(1600);
CN_in_sig(1818)	<=	VN_out_sig(1601);
CN_in_sig(3402)	<=	VN_out_sig(1602);
CN_in_sig(4458)	<=	VN_out_sig(1603);
CN_in_sig(962)	<=	VN_out_sig(1604);
CN_in_sig(1826)	<=	VN_out_sig(1605);
CN_in_sig(3410)	<=	VN_out_sig(1606);
CN_in_sig(4466)	<=	VN_out_sig(1607);
CN_in_sig(970)	<=	VN_out_sig(1608);
CN_in_sig(1834)	<=	VN_out_sig(1609);
CN_in_sig(3418)	<=	VN_out_sig(1610);
CN_in_sig(4474)	<=	VN_out_sig(1611);
CN_in_sig(978)	<=	VN_out_sig(1612);
CN_in_sig(1842)	<=	VN_out_sig(1613);
CN_in_sig(3426)	<=	VN_out_sig(1614);
CN_in_sig(4482)	<=	VN_out_sig(1615);
CN_in_sig(986)	<=	VN_out_sig(1616);
CN_in_sig(1850)	<=	VN_out_sig(1617);
CN_in_sig(3434)	<=	VN_out_sig(1618);
CN_in_sig(4490)	<=	VN_out_sig(1619);
CN_in_sig(994)	<=	VN_out_sig(1620);
CN_in_sig(1858)	<=	VN_out_sig(1621);
CN_in_sig(3442)	<=	VN_out_sig(1622);
CN_in_sig(4498)	<=	VN_out_sig(1623);
CN_in_sig(1002)	<=	VN_out_sig(1624);
CN_in_sig(1866)	<=	VN_out_sig(1625);
CN_in_sig(3450)	<=	VN_out_sig(1626);
CN_in_sig(4506)	<=	VN_out_sig(1627);
CN_in_sig(1010)	<=	VN_out_sig(1628);
CN_in_sig(1874)	<=	VN_out_sig(1629);
CN_in_sig(3026)	<=	VN_out_sig(1630);
CN_in_sig(4514)	<=	VN_out_sig(1631);
CN_in_sig(1018)	<=	VN_out_sig(1632);
CN_in_sig(1882)	<=	VN_out_sig(1633);
CN_in_sig(3034)	<=	VN_out_sig(1634);
CN_in_sig(4522)	<=	VN_out_sig(1635);
CN_in_sig(1026)	<=	VN_out_sig(1636);
CN_in_sig(1890)	<=	VN_out_sig(1637);
CN_in_sig(3042)	<=	VN_out_sig(1638);
CN_in_sig(4530)	<=	VN_out_sig(1639);
CN_in_sig(1034)	<=	VN_out_sig(1640);
CN_in_sig(1898)	<=	VN_out_sig(1641);
CN_in_sig(3050)	<=	VN_out_sig(1642);
CN_in_sig(4538)	<=	VN_out_sig(1643);
CN_in_sig(1042)	<=	VN_out_sig(1644);
CN_in_sig(1906)	<=	VN_out_sig(1645);
CN_in_sig(3058)	<=	VN_out_sig(1646);
CN_in_sig(4546)	<=	VN_out_sig(1647);
CN_in_sig(1050)	<=	VN_out_sig(1648);
CN_in_sig(1914)	<=	VN_out_sig(1649);
CN_in_sig(3066)	<=	VN_out_sig(1650);
CN_in_sig(4554)	<=	VN_out_sig(1651);
CN_in_sig(1058)	<=	VN_out_sig(1652);
CN_in_sig(1922)	<=	VN_out_sig(1653);
CN_in_sig(3074)	<=	VN_out_sig(1654);
CN_in_sig(4562)	<=	VN_out_sig(1655);
CN_in_sig(1066)	<=	VN_out_sig(1656);
CN_in_sig(1930)	<=	VN_out_sig(1657);
CN_in_sig(3082)	<=	VN_out_sig(1658);
CN_in_sig(4570)	<=	VN_out_sig(1659);
CN_in_sig(1074)	<=	VN_out_sig(1660);
CN_in_sig(1938)	<=	VN_out_sig(1661);
CN_in_sig(3090)	<=	VN_out_sig(1662);
CN_in_sig(4578)	<=	VN_out_sig(1663);
CN_in_sig(1082)	<=	VN_out_sig(1664);
CN_in_sig(1946)	<=	VN_out_sig(1665);
CN_in_sig(3098)	<=	VN_out_sig(1666);
CN_in_sig(4586)	<=	VN_out_sig(1667);
CN_in_sig(1090)	<=	VN_out_sig(1668);
CN_in_sig(1954)	<=	VN_out_sig(1669);
CN_in_sig(3106)	<=	VN_out_sig(1670);
CN_in_sig(4594)	<=	VN_out_sig(1671);
CN_in_sig(1098)	<=	VN_out_sig(1672);
CN_in_sig(1962)	<=	VN_out_sig(1673);
CN_in_sig(3114)	<=	VN_out_sig(1674);
CN_in_sig(4602)	<=	VN_out_sig(1675);
CN_in_sig(1106)	<=	VN_out_sig(1676);
CN_in_sig(1970)	<=	VN_out_sig(1677);
CN_in_sig(3122)	<=	VN_out_sig(1678);
CN_in_sig(4610)	<=	VN_out_sig(1679);
CN_in_sig(1114)	<=	VN_out_sig(1680);
CN_in_sig(1978)	<=	VN_out_sig(1681);
CN_in_sig(3130)	<=	VN_out_sig(1682);
CN_in_sig(4618)	<=	VN_out_sig(1683);
CN_in_sig(1122)	<=	VN_out_sig(1684);
CN_in_sig(1986)	<=	VN_out_sig(1685);
CN_in_sig(3138)	<=	VN_out_sig(1686);
CN_in_sig(4626)	<=	VN_out_sig(1687);
CN_in_sig(1130)	<=	VN_out_sig(1688);
CN_in_sig(1994)	<=	VN_out_sig(1689);
CN_in_sig(3146)	<=	VN_out_sig(1690);
CN_in_sig(4634)	<=	VN_out_sig(1691);
CN_in_sig(1138)	<=	VN_out_sig(1692);
CN_in_sig(2002)	<=	VN_out_sig(1693);
CN_in_sig(3154)	<=	VN_out_sig(1694);
CN_in_sig(4642)	<=	VN_out_sig(1695);
CN_in_sig(1146)	<=	VN_out_sig(1696);
CN_in_sig(2010)	<=	VN_out_sig(1697);
CN_in_sig(3162)	<=	VN_out_sig(1698);
CN_in_sig(4650)	<=	VN_out_sig(1699);
CN_in_sig(1154)	<=	VN_out_sig(1700);
CN_in_sig(2018)	<=	VN_out_sig(1701);
CN_in_sig(3170)	<=	VN_out_sig(1702);
CN_in_sig(4658)	<=	VN_out_sig(1703);
CN_in_sig(1162)	<=	VN_out_sig(1704);
CN_in_sig(2026)	<=	VN_out_sig(1705);
CN_in_sig(3178)	<=	VN_out_sig(1706);
CN_in_sig(4666)	<=	VN_out_sig(1707);
CN_in_sig(1170)	<=	VN_out_sig(1708);
CN_in_sig(2034)	<=	VN_out_sig(1709);
CN_in_sig(3186)	<=	VN_out_sig(1710);
CN_in_sig(4674)	<=	VN_out_sig(1711);
CN_in_sig(1178)	<=	VN_out_sig(1712);
CN_in_sig(2042)	<=	VN_out_sig(1713);
CN_in_sig(3194)	<=	VN_out_sig(1714);
CN_in_sig(4682)	<=	VN_out_sig(1715);
CN_in_sig(1186)	<=	VN_out_sig(1716);
CN_in_sig(2050)	<=	VN_out_sig(1717);
CN_in_sig(3202)	<=	VN_out_sig(1718);
CN_in_sig(4690)	<=	VN_out_sig(1719);
CN_in_sig(1194)	<=	VN_out_sig(1720);
CN_in_sig(2058)	<=	VN_out_sig(1721);
CN_in_sig(3210)	<=	VN_out_sig(1722);
CN_in_sig(4698)	<=	VN_out_sig(1723);
CN_in_sig(1202)	<=	VN_out_sig(1724);
CN_in_sig(2066)	<=	VN_out_sig(1725);
CN_in_sig(3218)	<=	VN_out_sig(1726);
CN_in_sig(4706)	<=	VN_out_sig(1727);
CN_in_sig(170)	<=	VN_out_sig(1728);
CN_in_sig(2514)	<=	VN_out_sig(1729);
CN_in_sig(2778)	<=	VN_out_sig(1730);
CN_in_sig(4114)	<=	VN_out_sig(1731);
CN_in_sig(178)	<=	VN_out_sig(1732);
CN_in_sig(2522)	<=	VN_out_sig(1733);
CN_in_sig(2786)	<=	VN_out_sig(1734);
CN_in_sig(4122)	<=	VN_out_sig(1735);
CN_in_sig(186)	<=	VN_out_sig(1736);
CN_in_sig(2530)	<=	VN_out_sig(1737);
CN_in_sig(2794)	<=	VN_out_sig(1738);
CN_in_sig(4130)	<=	VN_out_sig(1739);
CN_in_sig(194)	<=	VN_out_sig(1740);
CN_in_sig(2538)	<=	VN_out_sig(1741);
CN_in_sig(2802)	<=	VN_out_sig(1742);
CN_in_sig(4138)	<=	VN_out_sig(1743);
CN_in_sig(202)	<=	VN_out_sig(1744);
CN_in_sig(2546)	<=	VN_out_sig(1745);
CN_in_sig(2810)	<=	VN_out_sig(1746);
CN_in_sig(4146)	<=	VN_out_sig(1747);
CN_in_sig(210)	<=	VN_out_sig(1748);
CN_in_sig(2554)	<=	VN_out_sig(1749);
CN_in_sig(2818)	<=	VN_out_sig(1750);
CN_in_sig(4154)	<=	VN_out_sig(1751);
CN_in_sig(218)	<=	VN_out_sig(1752);
CN_in_sig(2562)	<=	VN_out_sig(1753);
CN_in_sig(2826)	<=	VN_out_sig(1754);
CN_in_sig(4162)	<=	VN_out_sig(1755);
CN_in_sig(226)	<=	VN_out_sig(1756);
CN_in_sig(2570)	<=	VN_out_sig(1757);
CN_in_sig(2834)	<=	VN_out_sig(1758);
CN_in_sig(4170)	<=	VN_out_sig(1759);
CN_in_sig(234)	<=	VN_out_sig(1760);
CN_in_sig(2578)	<=	VN_out_sig(1761);
CN_in_sig(2842)	<=	VN_out_sig(1762);
CN_in_sig(4178)	<=	VN_out_sig(1763);
CN_in_sig(242)	<=	VN_out_sig(1764);
CN_in_sig(2586)	<=	VN_out_sig(1765);
CN_in_sig(2850)	<=	VN_out_sig(1766);
CN_in_sig(4186)	<=	VN_out_sig(1767);
CN_in_sig(250)	<=	VN_out_sig(1768);
CN_in_sig(2162)	<=	VN_out_sig(1769);
CN_in_sig(2858)	<=	VN_out_sig(1770);
CN_in_sig(4194)	<=	VN_out_sig(1771);
CN_in_sig(258)	<=	VN_out_sig(1772);
CN_in_sig(2170)	<=	VN_out_sig(1773);
CN_in_sig(2866)	<=	VN_out_sig(1774);
CN_in_sig(4202)	<=	VN_out_sig(1775);
CN_in_sig(266)	<=	VN_out_sig(1776);
CN_in_sig(2178)	<=	VN_out_sig(1777);
CN_in_sig(2874)	<=	VN_out_sig(1778);
CN_in_sig(4210)	<=	VN_out_sig(1779);
CN_in_sig(274)	<=	VN_out_sig(1780);
CN_in_sig(2186)	<=	VN_out_sig(1781);
CN_in_sig(2882)	<=	VN_out_sig(1782);
CN_in_sig(4218)	<=	VN_out_sig(1783);
CN_in_sig(282)	<=	VN_out_sig(1784);
CN_in_sig(2194)	<=	VN_out_sig(1785);
CN_in_sig(2890)	<=	VN_out_sig(1786);
CN_in_sig(4226)	<=	VN_out_sig(1787);
CN_in_sig(290)	<=	VN_out_sig(1788);
CN_in_sig(2202)	<=	VN_out_sig(1789);
CN_in_sig(2898)	<=	VN_out_sig(1790);
CN_in_sig(4234)	<=	VN_out_sig(1791);
CN_in_sig(298)	<=	VN_out_sig(1792);
CN_in_sig(2210)	<=	VN_out_sig(1793);
CN_in_sig(2906)	<=	VN_out_sig(1794);
CN_in_sig(4242)	<=	VN_out_sig(1795);
CN_in_sig(306)	<=	VN_out_sig(1796);
CN_in_sig(2218)	<=	VN_out_sig(1797);
CN_in_sig(2914)	<=	VN_out_sig(1798);
CN_in_sig(4250)	<=	VN_out_sig(1799);
CN_in_sig(314)	<=	VN_out_sig(1800);
CN_in_sig(2226)	<=	VN_out_sig(1801);
CN_in_sig(2922)	<=	VN_out_sig(1802);
CN_in_sig(4258)	<=	VN_out_sig(1803);
CN_in_sig(322)	<=	VN_out_sig(1804);
CN_in_sig(2234)	<=	VN_out_sig(1805);
CN_in_sig(2930)	<=	VN_out_sig(1806);
CN_in_sig(4266)	<=	VN_out_sig(1807);
CN_in_sig(330)	<=	VN_out_sig(1808);
CN_in_sig(2242)	<=	VN_out_sig(1809);
CN_in_sig(2938)	<=	VN_out_sig(1810);
CN_in_sig(4274)	<=	VN_out_sig(1811);
CN_in_sig(338)	<=	VN_out_sig(1812);
CN_in_sig(2250)	<=	VN_out_sig(1813);
CN_in_sig(2946)	<=	VN_out_sig(1814);
CN_in_sig(4282)	<=	VN_out_sig(1815);
CN_in_sig(346)	<=	VN_out_sig(1816);
CN_in_sig(2258)	<=	VN_out_sig(1817);
CN_in_sig(2954)	<=	VN_out_sig(1818);
CN_in_sig(4290)	<=	VN_out_sig(1819);
CN_in_sig(354)	<=	VN_out_sig(1820);
CN_in_sig(2266)	<=	VN_out_sig(1821);
CN_in_sig(2962)	<=	VN_out_sig(1822);
CN_in_sig(4298)	<=	VN_out_sig(1823);
CN_in_sig(362)	<=	VN_out_sig(1824);
CN_in_sig(2274)	<=	VN_out_sig(1825);
CN_in_sig(2970)	<=	VN_out_sig(1826);
CN_in_sig(4306)	<=	VN_out_sig(1827);
CN_in_sig(370)	<=	VN_out_sig(1828);
CN_in_sig(2282)	<=	VN_out_sig(1829);
CN_in_sig(2978)	<=	VN_out_sig(1830);
CN_in_sig(4314)	<=	VN_out_sig(1831);
CN_in_sig(378)	<=	VN_out_sig(1832);
CN_in_sig(2290)	<=	VN_out_sig(1833);
CN_in_sig(2986)	<=	VN_out_sig(1834);
CN_in_sig(3890)	<=	VN_out_sig(1835);
CN_in_sig(386)	<=	VN_out_sig(1836);
CN_in_sig(2298)	<=	VN_out_sig(1837);
CN_in_sig(2994)	<=	VN_out_sig(1838);
CN_in_sig(3898)	<=	VN_out_sig(1839);
CN_in_sig(394)	<=	VN_out_sig(1840);
CN_in_sig(2306)	<=	VN_out_sig(1841);
CN_in_sig(3002)	<=	VN_out_sig(1842);
CN_in_sig(3906)	<=	VN_out_sig(1843);
CN_in_sig(402)	<=	VN_out_sig(1844);
CN_in_sig(2314)	<=	VN_out_sig(1845);
CN_in_sig(3010)	<=	VN_out_sig(1846);
CN_in_sig(3914)	<=	VN_out_sig(1847);
CN_in_sig(410)	<=	VN_out_sig(1848);
CN_in_sig(2322)	<=	VN_out_sig(1849);
CN_in_sig(3018)	<=	VN_out_sig(1850);
CN_in_sig(3922)	<=	VN_out_sig(1851);
CN_in_sig(418)	<=	VN_out_sig(1852);
CN_in_sig(2330)	<=	VN_out_sig(1853);
CN_in_sig(2594)	<=	VN_out_sig(1854);
CN_in_sig(3930)	<=	VN_out_sig(1855);
CN_in_sig(426)	<=	VN_out_sig(1856);
CN_in_sig(2338)	<=	VN_out_sig(1857);
CN_in_sig(2602)	<=	VN_out_sig(1858);
CN_in_sig(3938)	<=	VN_out_sig(1859);
CN_in_sig(2)	<=	VN_out_sig(1860);
CN_in_sig(2346)	<=	VN_out_sig(1861);
CN_in_sig(2610)	<=	VN_out_sig(1862);
CN_in_sig(3946)	<=	VN_out_sig(1863);
CN_in_sig(10)	<=	VN_out_sig(1864);
CN_in_sig(2354)	<=	VN_out_sig(1865);
CN_in_sig(2618)	<=	VN_out_sig(1866);
CN_in_sig(3954)	<=	VN_out_sig(1867);
CN_in_sig(18)	<=	VN_out_sig(1868);
CN_in_sig(2362)	<=	VN_out_sig(1869);
CN_in_sig(2626)	<=	VN_out_sig(1870);
CN_in_sig(3962)	<=	VN_out_sig(1871);
CN_in_sig(26)	<=	VN_out_sig(1872);
CN_in_sig(2370)	<=	VN_out_sig(1873);
CN_in_sig(2634)	<=	VN_out_sig(1874);
CN_in_sig(3970)	<=	VN_out_sig(1875);
CN_in_sig(34)	<=	VN_out_sig(1876);
CN_in_sig(2378)	<=	VN_out_sig(1877);
CN_in_sig(2642)	<=	VN_out_sig(1878);
CN_in_sig(3978)	<=	VN_out_sig(1879);
CN_in_sig(42)	<=	VN_out_sig(1880);
CN_in_sig(2386)	<=	VN_out_sig(1881);
CN_in_sig(2650)	<=	VN_out_sig(1882);
CN_in_sig(3986)	<=	VN_out_sig(1883);
CN_in_sig(50)	<=	VN_out_sig(1884);
CN_in_sig(2394)	<=	VN_out_sig(1885);
CN_in_sig(2658)	<=	VN_out_sig(1886);
CN_in_sig(3994)	<=	VN_out_sig(1887);
CN_in_sig(58)	<=	VN_out_sig(1888);
CN_in_sig(2402)	<=	VN_out_sig(1889);
CN_in_sig(2666)	<=	VN_out_sig(1890);
CN_in_sig(4002)	<=	VN_out_sig(1891);
CN_in_sig(66)	<=	VN_out_sig(1892);
CN_in_sig(2410)	<=	VN_out_sig(1893);
CN_in_sig(2674)	<=	VN_out_sig(1894);
CN_in_sig(4010)	<=	VN_out_sig(1895);
CN_in_sig(74)	<=	VN_out_sig(1896);
CN_in_sig(2418)	<=	VN_out_sig(1897);
CN_in_sig(2682)	<=	VN_out_sig(1898);
CN_in_sig(4018)	<=	VN_out_sig(1899);
CN_in_sig(82)	<=	VN_out_sig(1900);
CN_in_sig(2426)	<=	VN_out_sig(1901);
CN_in_sig(2690)	<=	VN_out_sig(1902);
CN_in_sig(4026)	<=	VN_out_sig(1903);
CN_in_sig(90)	<=	VN_out_sig(1904);
CN_in_sig(2434)	<=	VN_out_sig(1905);
CN_in_sig(2698)	<=	VN_out_sig(1906);
CN_in_sig(4034)	<=	VN_out_sig(1907);
CN_in_sig(98)	<=	VN_out_sig(1908);
CN_in_sig(2442)	<=	VN_out_sig(1909);
CN_in_sig(2706)	<=	VN_out_sig(1910);
CN_in_sig(4042)	<=	VN_out_sig(1911);
CN_in_sig(106)	<=	VN_out_sig(1912);
CN_in_sig(2450)	<=	VN_out_sig(1913);
CN_in_sig(2714)	<=	VN_out_sig(1914);
CN_in_sig(4050)	<=	VN_out_sig(1915);
CN_in_sig(114)	<=	VN_out_sig(1916);
CN_in_sig(2458)	<=	VN_out_sig(1917);
CN_in_sig(2722)	<=	VN_out_sig(1918);
CN_in_sig(4058)	<=	VN_out_sig(1919);
CN_in_sig(122)	<=	VN_out_sig(1920);
CN_in_sig(2466)	<=	VN_out_sig(1921);
CN_in_sig(2730)	<=	VN_out_sig(1922);
CN_in_sig(4066)	<=	VN_out_sig(1923);
CN_in_sig(130)	<=	VN_out_sig(1924);
CN_in_sig(2474)	<=	VN_out_sig(1925);
CN_in_sig(2738)	<=	VN_out_sig(1926);
CN_in_sig(4074)	<=	VN_out_sig(1927);
CN_in_sig(138)	<=	VN_out_sig(1928);
CN_in_sig(2482)	<=	VN_out_sig(1929);
CN_in_sig(2746)	<=	VN_out_sig(1930);
CN_in_sig(4082)	<=	VN_out_sig(1931);
CN_in_sig(146)	<=	VN_out_sig(1932);
CN_in_sig(2490)	<=	VN_out_sig(1933);
CN_in_sig(2754)	<=	VN_out_sig(1934);
CN_in_sig(4090)	<=	VN_out_sig(1935);
CN_in_sig(154)	<=	VN_out_sig(1936);
CN_in_sig(2498)	<=	VN_out_sig(1937);
CN_in_sig(2762)	<=	VN_out_sig(1938);
CN_in_sig(4098)	<=	VN_out_sig(1939);
CN_in_sig(162)	<=	VN_out_sig(1940);
CN_in_sig(2506)	<=	VN_out_sig(1941);
CN_in_sig(2770)	<=	VN_out_sig(1942);
CN_in_sig(4106)	<=	VN_out_sig(1943);
CN_in_sig(307)	<=	VN_out_sig(1944);
CN_in_sig(1571)	<=	VN_out_sig(1945);
CN_in_sig(2875)	<=	VN_out_sig(1946);
CN_in_sig(4915)	<=	VN_out_sig(1947);
CN_in_sig(315)	<=	VN_out_sig(1948);
CN_in_sig(1579)	<=	VN_out_sig(1949);
CN_in_sig(2883)	<=	VN_out_sig(1950);
CN_in_sig(4923)	<=	VN_out_sig(1951);
CN_in_sig(323)	<=	VN_out_sig(1952);
CN_in_sig(1587)	<=	VN_out_sig(1953);
CN_in_sig(2891)	<=	VN_out_sig(1954);
CN_in_sig(4931)	<=	VN_out_sig(1955);
CN_in_sig(331)	<=	VN_out_sig(1956);
CN_in_sig(1595)	<=	VN_out_sig(1957);
CN_in_sig(2899)	<=	VN_out_sig(1958);
CN_in_sig(4939)	<=	VN_out_sig(1959);
CN_in_sig(339)	<=	VN_out_sig(1960);
CN_in_sig(1603)	<=	VN_out_sig(1961);
CN_in_sig(2907)	<=	VN_out_sig(1962);
CN_in_sig(4947)	<=	VN_out_sig(1963);
CN_in_sig(347)	<=	VN_out_sig(1964);
CN_in_sig(1611)	<=	VN_out_sig(1965);
CN_in_sig(2915)	<=	VN_out_sig(1966);
CN_in_sig(4955)	<=	VN_out_sig(1967);
CN_in_sig(355)	<=	VN_out_sig(1968);
CN_in_sig(1619)	<=	VN_out_sig(1969);
CN_in_sig(2923)	<=	VN_out_sig(1970);
CN_in_sig(4963)	<=	VN_out_sig(1971);
CN_in_sig(363)	<=	VN_out_sig(1972);
CN_in_sig(1627)	<=	VN_out_sig(1973);
CN_in_sig(2931)	<=	VN_out_sig(1974);
CN_in_sig(4971)	<=	VN_out_sig(1975);
CN_in_sig(371)	<=	VN_out_sig(1976);
CN_in_sig(1635)	<=	VN_out_sig(1977);
CN_in_sig(2939)	<=	VN_out_sig(1978);
CN_in_sig(4979)	<=	VN_out_sig(1979);
CN_in_sig(379)	<=	VN_out_sig(1980);
CN_in_sig(1643)	<=	VN_out_sig(1981);
CN_in_sig(2947)	<=	VN_out_sig(1982);
CN_in_sig(4987)	<=	VN_out_sig(1983);
CN_in_sig(387)	<=	VN_out_sig(1984);
CN_in_sig(1651)	<=	VN_out_sig(1985);
CN_in_sig(2955)	<=	VN_out_sig(1986);
CN_in_sig(4995)	<=	VN_out_sig(1987);
CN_in_sig(395)	<=	VN_out_sig(1988);
CN_in_sig(1659)	<=	VN_out_sig(1989);
CN_in_sig(2963)	<=	VN_out_sig(1990);
CN_in_sig(5003)	<=	VN_out_sig(1991);
CN_in_sig(403)	<=	VN_out_sig(1992);
CN_in_sig(1667)	<=	VN_out_sig(1993);
CN_in_sig(2971)	<=	VN_out_sig(1994);
CN_in_sig(5011)	<=	VN_out_sig(1995);
CN_in_sig(411)	<=	VN_out_sig(1996);
CN_in_sig(1675)	<=	VN_out_sig(1997);
CN_in_sig(2979)	<=	VN_out_sig(1998);
CN_in_sig(5019)	<=	VN_out_sig(1999);
CN_in_sig(419)	<=	VN_out_sig(2000);
CN_in_sig(1683)	<=	VN_out_sig(2001);
CN_in_sig(2987)	<=	VN_out_sig(2002);
CN_in_sig(5027)	<=	VN_out_sig(2003);
CN_in_sig(427)	<=	VN_out_sig(2004);
CN_in_sig(1691)	<=	VN_out_sig(2005);
CN_in_sig(2995)	<=	VN_out_sig(2006);
CN_in_sig(5035)	<=	VN_out_sig(2007);
CN_in_sig(3)	<=	VN_out_sig(2008);
CN_in_sig(1699)	<=	VN_out_sig(2009);
CN_in_sig(3003)	<=	VN_out_sig(2010);
CN_in_sig(5043)	<=	VN_out_sig(2011);
CN_in_sig(11)	<=	VN_out_sig(2012);
CN_in_sig(1707)	<=	VN_out_sig(2013);
CN_in_sig(3011)	<=	VN_out_sig(2014);
CN_in_sig(5051)	<=	VN_out_sig(2015);
CN_in_sig(19)	<=	VN_out_sig(2016);
CN_in_sig(1715)	<=	VN_out_sig(2017);
CN_in_sig(3019)	<=	VN_out_sig(2018);
CN_in_sig(5059)	<=	VN_out_sig(2019);
CN_in_sig(27)	<=	VN_out_sig(2020);
CN_in_sig(1723)	<=	VN_out_sig(2021);
CN_in_sig(2595)	<=	VN_out_sig(2022);
CN_in_sig(5067)	<=	VN_out_sig(2023);
CN_in_sig(35)	<=	VN_out_sig(2024);
CN_in_sig(1299)	<=	VN_out_sig(2025);
CN_in_sig(2603)	<=	VN_out_sig(2026);
CN_in_sig(5075)	<=	VN_out_sig(2027);
CN_in_sig(43)	<=	VN_out_sig(2028);
CN_in_sig(1307)	<=	VN_out_sig(2029);
CN_in_sig(2611)	<=	VN_out_sig(2030);
CN_in_sig(5083)	<=	VN_out_sig(2031);
CN_in_sig(51)	<=	VN_out_sig(2032);
CN_in_sig(1315)	<=	VN_out_sig(2033);
CN_in_sig(2619)	<=	VN_out_sig(2034);
CN_in_sig(5091)	<=	VN_out_sig(2035);
CN_in_sig(59)	<=	VN_out_sig(2036);
CN_in_sig(1323)	<=	VN_out_sig(2037);
CN_in_sig(2627)	<=	VN_out_sig(2038);
CN_in_sig(5099)	<=	VN_out_sig(2039);
CN_in_sig(67)	<=	VN_out_sig(2040);
CN_in_sig(1331)	<=	VN_out_sig(2041);
CN_in_sig(2635)	<=	VN_out_sig(2042);
CN_in_sig(5107)	<=	VN_out_sig(2043);
CN_in_sig(75)	<=	VN_out_sig(2044);
CN_in_sig(1339)	<=	VN_out_sig(2045);
CN_in_sig(2643)	<=	VN_out_sig(2046);
CN_in_sig(5115)	<=	VN_out_sig(2047);
CN_in_sig(83)	<=	VN_out_sig(2048);
CN_in_sig(1347)	<=	VN_out_sig(2049);
CN_in_sig(2651)	<=	VN_out_sig(2050);
CN_in_sig(5123)	<=	VN_out_sig(2051);
CN_in_sig(91)	<=	VN_out_sig(2052);
CN_in_sig(1355)	<=	VN_out_sig(2053);
CN_in_sig(2659)	<=	VN_out_sig(2054);
CN_in_sig(5131)	<=	VN_out_sig(2055);
CN_in_sig(99)	<=	VN_out_sig(2056);
CN_in_sig(1363)	<=	VN_out_sig(2057);
CN_in_sig(2667)	<=	VN_out_sig(2058);
CN_in_sig(5139)	<=	VN_out_sig(2059);
CN_in_sig(107)	<=	VN_out_sig(2060);
CN_in_sig(1371)	<=	VN_out_sig(2061);
CN_in_sig(2675)	<=	VN_out_sig(2062);
CN_in_sig(5147)	<=	VN_out_sig(2063);
CN_in_sig(115)	<=	VN_out_sig(2064);
CN_in_sig(1379)	<=	VN_out_sig(2065);
CN_in_sig(2683)	<=	VN_out_sig(2066);
CN_in_sig(5155)	<=	VN_out_sig(2067);
CN_in_sig(123)	<=	VN_out_sig(2068);
CN_in_sig(1387)	<=	VN_out_sig(2069);
CN_in_sig(2691)	<=	VN_out_sig(2070);
CN_in_sig(5163)	<=	VN_out_sig(2071);
CN_in_sig(131)	<=	VN_out_sig(2072);
CN_in_sig(1395)	<=	VN_out_sig(2073);
CN_in_sig(2699)	<=	VN_out_sig(2074);
CN_in_sig(5171)	<=	VN_out_sig(2075);
CN_in_sig(139)	<=	VN_out_sig(2076);
CN_in_sig(1403)	<=	VN_out_sig(2077);
CN_in_sig(2707)	<=	VN_out_sig(2078);
CN_in_sig(5179)	<=	VN_out_sig(2079);
CN_in_sig(147)	<=	VN_out_sig(2080);
CN_in_sig(1411)	<=	VN_out_sig(2081);
CN_in_sig(2715)	<=	VN_out_sig(2082);
CN_in_sig(4755)	<=	VN_out_sig(2083);
CN_in_sig(155)	<=	VN_out_sig(2084);
CN_in_sig(1419)	<=	VN_out_sig(2085);
CN_in_sig(2723)	<=	VN_out_sig(2086);
CN_in_sig(4763)	<=	VN_out_sig(2087);
CN_in_sig(163)	<=	VN_out_sig(2088);
CN_in_sig(1427)	<=	VN_out_sig(2089);
CN_in_sig(2731)	<=	VN_out_sig(2090);
CN_in_sig(4771)	<=	VN_out_sig(2091);
CN_in_sig(171)	<=	VN_out_sig(2092);
CN_in_sig(1435)	<=	VN_out_sig(2093);
CN_in_sig(2739)	<=	VN_out_sig(2094);
CN_in_sig(4779)	<=	VN_out_sig(2095);
CN_in_sig(179)	<=	VN_out_sig(2096);
CN_in_sig(1443)	<=	VN_out_sig(2097);
CN_in_sig(2747)	<=	VN_out_sig(2098);
CN_in_sig(4787)	<=	VN_out_sig(2099);
CN_in_sig(187)	<=	VN_out_sig(2100);
CN_in_sig(1451)	<=	VN_out_sig(2101);
CN_in_sig(2755)	<=	VN_out_sig(2102);
CN_in_sig(4795)	<=	VN_out_sig(2103);
CN_in_sig(195)	<=	VN_out_sig(2104);
CN_in_sig(1459)	<=	VN_out_sig(2105);
CN_in_sig(2763)	<=	VN_out_sig(2106);
CN_in_sig(4803)	<=	VN_out_sig(2107);
CN_in_sig(203)	<=	VN_out_sig(2108);
CN_in_sig(1467)	<=	VN_out_sig(2109);
CN_in_sig(2771)	<=	VN_out_sig(2110);
CN_in_sig(4811)	<=	VN_out_sig(2111);
CN_in_sig(211)	<=	VN_out_sig(2112);
CN_in_sig(1475)	<=	VN_out_sig(2113);
CN_in_sig(2779)	<=	VN_out_sig(2114);
CN_in_sig(4819)	<=	VN_out_sig(2115);
CN_in_sig(219)	<=	VN_out_sig(2116);
CN_in_sig(1483)	<=	VN_out_sig(2117);
CN_in_sig(2787)	<=	VN_out_sig(2118);
CN_in_sig(4827)	<=	VN_out_sig(2119);
CN_in_sig(227)	<=	VN_out_sig(2120);
CN_in_sig(1491)	<=	VN_out_sig(2121);
CN_in_sig(2795)	<=	VN_out_sig(2122);
CN_in_sig(4835)	<=	VN_out_sig(2123);
CN_in_sig(235)	<=	VN_out_sig(2124);
CN_in_sig(1499)	<=	VN_out_sig(2125);
CN_in_sig(2803)	<=	VN_out_sig(2126);
CN_in_sig(4843)	<=	VN_out_sig(2127);
CN_in_sig(243)	<=	VN_out_sig(2128);
CN_in_sig(1507)	<=	VN_out_sig(2129);
CN_in_sig(2811)	<=	VN_out_sig(2130);
CN_in_sig(4851)	<=	VN_out_sig(2131);
CN_in_sig(251)	<=	VN_out_sig(2132);
CN_in_sig(1515)	<=	VN_out_sig(2133);
CN_in_sig(2819)	<=	VN_out_sig(2134);
CN_in_sig(4859)	<=	VN_out_sig(2135);
CN_in_sig(259)	<=	VN_out_sig(2136);
CN_in_sig(1523)	<=	VN_out_sig(2137);
CN_in_sig(2827)	<=	VN_out_sig(2138);
CN_in_sig(4867)	<=	VN_out_sig(2139);
CN_in_sig(267)	<=	VN_out_sig(2140);
CN_in_sig(1531)	<=	VN_out_sig(2141);
CN_in_sig(2835)	<=	VN_out_sig(2142);
CN_in_sig(4875)	<=	VN_out_sig(2143);
CN_in_sig(275)	<=	VN_out_sig(2144);
CN_in_sig(1539)	<=	VN_out_sig(2145);
CN_in_sig(2843)	<=	VN_out_sig(2146);
CN_in_sig(4883)	<=	VN_out_sig(2147);
CN_in_sig(283)	<=	VN_out_sig(2148);
CN_in_sig(1547)	<=	VN_out_sig(2149);
CN_in_sig(2851)	<=	VN_out_sig(2150);
CN_in_sig(4891)	<=	VN_out_sig(2151);
CN_in_sig(291)	<=	VN_out_sig(2152);
CN_in_sig(1555)	<=	VN_out_sig(2153);
CN_in_sig(2859)	<=	VN_out_sig(2154);
CN_in_sig(4899)	<=	VN_out_sig(2155);
CN_in_sig(299)	<=	VN_out_sig(2156);
CN_in_sig(1563)	<=	VN_out_sig(2157);
CN_in_sig(2867)	<=	VN_out_sig(2158);
CN_in_sig(4907)	<=	VN_out_sig(2159);
CN_in_sig(635)	<=	VN_out_sig(2160);
CN_in_sig(2451)	<=	VN_out_sig(2161);
CN_in_sig(3419)	<=	VN_out_sig(2162);
CN_in_sig(4299)	<=	VN_out_sig(2163);
CN_in_sig(643)	<=	VN_out_sig(2164);
CN_in_sig(2459)	<=	VN_out_sig(2165);
CN_in_sig(3427)	<=	VN_out_sig(2166);
CN_in_sig(4307)	<=	VN_out_sig(2167);
CN_in_sig(651)	<=	VN_out_sig(2168);
CN_in_sig(2467)	<=	VN_out_sig(2169);
CN_in_sig(3435)	<=	VN_out_sig(2170);
CN_in_sig(4315)	<=	VN_out_sig(2171);
CN_in_sig(659)	<=	VN_out_sig(2172);
CN_in_sig(2475)	<=	VN_out_sig(2173);
CN_in_sig(3443)	<=	VN_out_sig(2174);
CN_in_sig(3891)	<=	VN_out_sig(2175);
CN_in_sig(667)	<=	VN_out_sig(2176);
CN_in_sig(2483)	<=	VN_out_sig(2177);
CN_in_sig(3451)	<=	VN_out_sig(2178);
CN_in_sig(3899)	<=	VN_out_sig(2179);
CN_in_sig(675)	<=	VN_out_sig(2180);
CN_in_sig(2491)	<=	VN_out_sig(2181);
CN_in_sig(3027)	<=	VN_out_sig(2182);
CN_in_sig(3907)	<=	VN_out_sig(2183);
CN_in_sig(683)	<=	VN_out_sig(2184);
CN_in_sig(2499)	<=	VN_out_sig(2185);
CN_in_sig(3035)	<=	VN_out_sig(2186);
CN_in_sig(3915)	<=	VN_out_sig(2187);
CN_in_sig(691)	<=	VN_out_sig(2188);
CN_in_sig(2507)	<=	VN_out_sig(2189);
CN_in_sig(3043)	<=	VN_out_sig(2190);
CN_in_sig(3923)	<=	VN_out_sig(2191);
CN_in_sig(699)	<=	VN_out_sig(2192);
CN_in_sig(2515)	<=	VN_out_sig(2193);
CN_in_sig(3051)	<=	VN_out_sig(2194);
CN_in_sig(3931)	<=	VN_out_sig(2195);
CN_in_sig(707)	<=	VN_out_sig(2196);
CN_in_sig(2523)	<=	VN_out_sig(2197);
CN_in_sig(3059)	<=	VN_out_sig(2198);
CN_in_sig(3939)	<=	VN_out_sig(2199);
CN_in_sig(715)	<=	VN_out_sig(2200);
CN_in_sig(2531)	<=	VN_out_sig(2201);
CN_in_sig(3067)	<=	VN_out_sig(2202);
CN_in_sig(3947)	<=	VN_out_sig(2203);
CN_in_sig(723)	<=	VN_out_sig(2204);
CN_in_sig(2539)	<=	VN_out_sig(2205);
CN_in_sig(3075)	<=	VN_out_sig(2206);
CN_in_sig(3955)	<=	VN_out_sig(2207);
CN_in_sig(731)	<=	VN_out_sig(2208);
CN_in_sig(2547)	<=	VN_out_sig(2209);
CN_in_sig(3083)	<=	VN_out_sig(2210);
CN_in_sig(3963)	<=	VN_out_sig(2211);
CN_in_sig(739)	<=	VN_out_sig(2212);
CN_in_sig(2555)	<=	VN_out_sig(2213);
CN_in_sig(3091)	<=	VN_out_sig(2214);
CN_in_sig(3971)	<=	VN_out_sig(2215);
CN_in_sig(747)	<=	VN_out_sig(2216);
CN_in_sig(2563)	<=	VN_out_sig(2217);
CN_in_sig(3099)	<=	VN_out_sig(2218);
CN_in_sig(3979)	<=	VN_out_sig(2219);
CN_in_sig(755)	<=	VN_out_sig(2220);
CN_in_sig(2571)	<=	VN_out_sig(2221);
CN_in_sig(3107)	<=	VN_out_sig(2222);
CN_in_sig(3987)	<=	VN_out_sig(2223);
CN_in_sig(763)	<=	VN_out_sig(2224);
CN_in_sig(2579)	<=	VN_out_sig(2225);
CN_in_sig(3115)	<=	VN_out_sig(2226);
CN_in_sig(3995)	<=	VN_out_sig(2227);
CN_in_sig(771)	<=	VN_out_sig(2228);
CN_in_sig(2587)	<=	VN_out_sig(2229);
CN_in_sig(3123)	<=	VN_out_sig(2230);
CN_in_sig(4003)	<=	VN_out_sig(2231);
CN_in_sig(779)	<=	VN_out_sig(2232);
CN_in_sig(2163)	<=	VN_out_sig(2233);
CN_in_sig(3131)	<=	VN_out_sig(2234);
CN_in_sig(4011)	<=	VN_out_sig(2235);
CN_in_sig(787)	<=	VN_out_sig(2236);
CN_in_sig(2171)	<=	VN_out_sig(2237);
CN_in_sig(3139)	<=	VN_out_sig(2238);
CN_in_sig(4019)	<=	VN_out_sig(2239);
CN_in_sig(795)	<=	VN_out_sig(2240);
CN_in_sig(2179)	<=	VN_out_sig(2241);
CN_in_sig(3147)	<=	VN_out_sig(2242);
CN_in_sig(4027)	<=	VN_out_sig(2243);
CN_in_sig(803)	<=	VN_out_sig(2244);
CN_in_sig(2187)	<=	VN_out_sig(2245);
CN_in_sig(3155)	<=	VN_out_sig(2246);
CN_in_sig(4035)	<=	VN_out_sig(2247);
CN_in_sig(811)	<=	VN_out_sig(2248);
CN_in_sig(2195)	<=	VN_out_sig(2249);
CN_in_sig(3163)	<=	VN_out_sig(2250);
CN_in_sig(4043)	<=	VN_out_sig(2251);
CN_in_sig(819)	<=	VN_out_sig(2252);
CN_in_sig(2203)	<=	VN_out_sig(2253);
CN_in_sig(3171)	<=	VN_out_sig(2254);
CN_in_sig(4051)	<=	VN_out_sig(2255);
CN_in_sig(827)	<=	VN_out_sig(2256);
CN_in_sig(2211)	<=	VN_out_sig(2257);
CN_in_sig(3179)	<=	VN_out_sig(2258);
CN_in_sig(4059)	<=	VN_out_sig(2259);
CN_in_sig(835)	<=	VN_out_sig(2260);
CN_in_sig(2219)	<=	VN_out_sig(2261);
CN_in_sig(3187)	<=	VN_out_sig(2262);
CN_in_sig(4067)	<=	VN_out_sig(2263);
CN_in_sig(843)	<=	VN_out_sig(2264);
CN_in_sig(2227)	<=	VN_out_sig(2265);
CN_in_sig(3195)	<=	VN_out_sig(2266);
CN_in_sig(4075)	<=	VN_out_sig(2267);
CN_in_sig(851)	<=	VN_out_sig(2268);
CN_in_sig(2235)	<=	VN_out_sig(2269);
CN_in_sig(3203)	<=	VN_out_sig(2270);
CN_in_sig(4083)	<=	VN_out_sig(2271);
CN_in_sig(859)	<=	VN_out_sig(2272);
CN_in_sig(2243)	<=	VN_out_sig(2273);
CN_in_sig(3211)	<=	VN_out_sig(2274);
CN_in_sig(4091)	<=	VN_out_sig(2275);
CN_in_sig(435)	<=	VN_out_sig(2276);
CN_in_sig(2251)	<=	VN_out_sig(2277);
CN_in_sig(3219)	<=	VN_out_sig(2278);
CN_in_sig(4099)	<=	VN_out_sig(2279);
CN_in_sig(443)	<=	VN_out_sig(2280);
CN_in_sig(2259)	<=	VN_out_sig(2281);
CN_in_sig(3227)	<=	VN_out_sig(2282);
CN_in_sig(4107)	<=	VN_out_sig(2283);
CN_in_sig(451)	<=	VN_out_sig(2284);
CN_in_sig(2267)	<=	VN_out_sig(2285);
CN_in_sig(3235)	<=	VN_out_sig(2286);
CN_in_sig(4115)	<=	VN_out_sig(2287);
CN_in_sig(459)	<=	VN_out_sig(2288);
CN_in_sig(2275)	<=	VN_out_sig(2289);
CN_in_sig(3243)	<=	VN_out_sig(2290);
CN_in_sig(4123)	<=	VN_out_sig(2291);
CN_in_sig(467)	<=	VN_out_sig(2292);
CN_in_sig(2283)	<=	VN_out_sig(2293);
CN_in_sig(3251)	<=	VN_out_sig(2294);
CN_in_sig(4131)	<=	VN_out_sig(2295);
CN_in_sig(475)	<=	VN_out_sig(2296);
CN_in_sig(2291)	<=	VN_out_sig(2297);
CN_in_sig(3259)	<=	VN_out_sig(2298);
CN_in_sig(4139)	<=	VN_out_sig(2299);
CN_in_sig(483)	<=	VN_out_sig(2300);
CN_in_sig(2299)	<=	VN_out_sig(2301);
CN_in_sig(3267)	<=	VN_out_sig(2302);
CN_in_sig(4147)	<=	VN_out_sig(2303);
CN_in_sig(491)	<=	VN_out_sig(2304);
CN_in_sig(2307)	<=	VN_out_sig(2305);
CN_in_sig(3275)	<=	VN_out_sig(2306);
CN_in_sig(4155)	<=	VN_out_sig(2307);
CN_in_sig(499)	<=	VN_out_sig(2308);
CN_in_sig(2315)	<=	VN_out_sig(2309);
CN_in_sig(3283)	<=	VN_out_sig(2310);
CN_in_sig(4163)	<=	VN_out_sig(2311);
CN_in_sig(507)	<=	VN_out_sig(2312);
CN_in_sig(2323)	<=	VN_out_sig(2313);
CN_in_sig(3291)	<=	VN_out_sig(2314);
CN_in_sig(4171)	<=	VN_out_sig(2315);
CN_in_sig(515)	<=	VN_out_sig(2316);
CN_in_sig(2331)	<=	VN_out_sig(2317);
CN_in_sig(3299)	<=	VN_out_sig(2318);
CN_in_sig(4179)	<=	VN_out_sig(2319);
CN_in_sig(523)	<=	VN_out_sig(2320);
CN_in_sig(2339)	<=	VN_out_sig(2321);
CN_in_sig(3307)	<=	VN_out_sig(2322);
CN_in_sig(4187)	<=	VN_out_sig(2323);
CN_in_sig(531)	<=	VN_out_sig(2324);
CN_in_sig(2347)	<=	VN_out_sig(2325);
CN_in_sig(3315)	<=	VN_out_sig(2326);
CN_in_sig(4195)	<=	VN_out_sig(2327);
CN_in_sig(539)	<=	VN_out_sig(2328);
CN_in_sig(2355)	<=	VN_out_sig(2329);
CN_in_sig(3323)	<=	VN_out_sig(2330);
CN_in_sig(4203)	<=	VN_out_sig(2331);
CN_in_sig(547)	<=	VN_out_sig(2332);
CN_in_sig(2363)	<=	VN_out_sig(2333);
CN_in_sig(3331)	<=	VN_out_sig(2334);
CN_in_sig(4211)	<=	VN_out_sig(2335);
CN_in_sig(555)	<=	VN_out_sig(2336);
CN_in_sig(2371)	<=	VN_out_sig(2337);
CN_in_sig(3339)	<=	VN_out_sig(2338);
CN_in_sig(4219)	<=	VN_out_sig(2339);
CN_in_sig(563)	<=	VN_out_sig(2340);
CN_in_sig(2379)	<=	VN_out_sig(2341);
CN_in_sig(3347)	<=	VN_out_sig(2342);
CN_in_sig(4227)	<=	VN_out_sig(2343);
CN_in_sig(571)	<=	VN_out_sig(2344);
CN_in_sig(2387)	<=	VN_out_sig(2345);
CN_in_sig(3355)	<=	VN_out_sig(2346);
CN_in_sig(4235)	<=	VN_out_sig(2347);
CN_in_sig(579)	<=	VN_out_sig(2348);
CN_in_sig(2395)	<=	VN_out_sig(2349);
CN_in_sig(3363)	<=	VN_out_sig(2350);
CN_in_sig(4243)	<=	VN_out_sig(2351);
CN_in_sig(587)	<=	VN_out_sig(2352);
CN_in_sig(2403)	<=	VN_out_sig(2353);
CN_in_sig(3371)	<=	VN_out_sig(2354);
CN_in_sig(4251)	<=	VN_out_sig(2355);
CN_in_sig(595)	<=	VN_out_sig(2356);
CN_in_sig(2411)	<=	VN_out_sig(2357);
CN_in_sig(3379)	<=	VN_out_sig(2358);
CN_in_sig(4259)	<=	VN_out_sig(2359);
CN_in_sig(603)	<=	VN_out_sig(2360);
CN_in_sig(2419)	<=	VN_out_sig(2361);
CN_in_sig(3387)	<=	VN_out_sig(2362);
CN_in_sig(4267)	<=	VN_out_sig(2363);
CN_in_sig(611)	<=	VN_out_sig(2364);
CN_in_sig(2427)	<=	VN_out_sig(2365);
CN_in_sig(3395)	<=	VN_out_sig(2366);
CN_in_sig(4275)	<=	VN_out_sig(2367);
CN_in_sig(619)	<=	VN_out_sig(2368);
CN_in_sig(2435)	<=	VN_out_sig(2369);
CN_in_sig(3403)	<=	VN_out_sig(2370);
CN_in_sig(4283)	<=	VN_out_sig(2371);
CN_in_sig(627)	<=	VN_out_sig(2372);
CN_in_sig(2443)	<=	VN_out_sig(2373);
CN_in_sig(3411)	<=	VN_out_sig(2374);
CN_in_sig(4291)	<=	VN_out_sig(2375);
CN_in_sig(1283)	<=	VN_out_sig(2376);
CN_in_sig(1811)	<=	VN_out_sig(2377);
CN_in_sig(3883)	<=	VN_out_sig(2378);
CN_in_sig(4651)	<=	VN_out_sig(2379);
CN_in_sig(1291)	<=	VN_out_sig(2380);
CN_in_sig(1819)	<=	VN_out_sig(2381);
CN_in_sig(3459)	<=	VN_out_sig(2382);
CN_in_sig(4659)	<=	VN_out_sig(2383);
CN_in_sig(867)	<=	VN_out_sig(2384);
CN_in_sig(1827)	<=	VN_out_sig(2385);
CN_in_sig(3467)	<=	VN_out_sig(2386);
CN_in_sig(4667)	<=	VN_out_sig(2387);
CN_in_sig(875)	<=	VN_out_sig(2388);
CN_in_sig(1835)	<=	VN_out_sig(2389);
CN_in_sig(3475)	<=	VN_out_sig(2390);
CN_in_sig(4675)	<=	VN_out_sig(2391);
CN_in_sig(883)	<=	VN_out_sig(2392);
CN_in_sig(1843)	<=	VN_out_sig(2393);
CN_in_sig(3483)	<=	VN_out_sig(2394);
CN_in_sig(4683)	<=	VN_out_sig(2395);
CN_in_sig(891)	<=	VN_out_sig(2396);
CN_in_sig(1851)	<=	VN_out_sig(2397);
CN_in_sig(3491)	<=	VN_out_sig(2398);
CN_in_sig(4691)	<=	VN_out_sig(2399);
CN_in_sig(899)	<=	VN_out_sig(2400);
CN_in_sig(1859)	<=	VN_out_sig(2401);
CN_in_sig(3499)	<=	VN_out_sig(2402);
CN_in_sig(4699)	<=	VN_out_sig(2403);
CN_in_sig(907)	<=	VN_out_sig(2404);
CN_in_sig(1867)	<=	VN_out_sig(2405);
CN_in_sig(3507)	<=	VN_out_sig(2406);
CN_in_sig(4707)	<=	VN_out_sig(2407);
CN_in_sig(915)	<=	VN_out_sig(2408);
CN_in_sig(1875)	<=	VN_out_sig(2409);
CN_in_sig(3515)	<=	VN_out_sig(2410);
CN_in_sig(4715)	<=	VN_out_sig(2411);
CN_in_sig(923)	<=	VN_out_sig(2412);
CN_in_sig(1883)	<=	VN_out_sig(2413);
CN_in_sig(3523)	<=	VN_out_sig(2414);
CN_in_sig(4723)	<=	VN_out_sig(2415);
CN_in_sig(931)	<=	VN_out_sig(2416);
CN_in_sig(1891)	<=	VN_out_sig(2417);
CN_in_sig(3531)	<=	VN_out_sig(2418);
CN_in_sig(4731)	<=	VN_out_sig(2419);
CN_in_sig(939)	<=	VN_out_sig(2420);
CN_in_sig(1899)	<=	VN_out_sig(2421);
CN_in_sig(3539)	<=	VN_out_sig(2422);
CN_in_sig(4739)	<=	VN_out_sig(2423);
CN_in_sig(947)	<=	VN_out_sig(2424);
CN_in_sig(1907)	<=	VN_out_sig(2425);
CN_in_sig(3547)	<=	VN_out_sig(2426);
CN_in_sig(4747)	<=	VN_out_sig(2427);
CN_in_sig(955)	<=	VN_out_sig(2428);
CN_in_sig(1915)	<=	VN_out_sig(2429);
CN_in_sig(3555)	<=	VN_out_sig(2430);
CN_in_sig(4323)	<=	VN_out_sig(2431);
CN_in_sig(963)	<=	VN_out_sig(2432);
CN_in_sig(1923)	<=	VN_out_sig(2433);
CN_in_sig(3563)	<=	VN_out_sig(2434);
CN_in_sig(4331)	<=	VN_out_sig(2435);
CN_in_sig(971)	<=	VN_out_sig(2436);
CN_in_sig(1931)	<=	VN_out_sig(2437);
CN_in_sig(3571)	<=	VN_out_sig(2438);
CN_in_sig(4339)	<=	VN_out_sig(2439);
CN_in_sig(979)	<=	VN_out_sig(2440);
CN_in_sig(1939)	<=	VN_out_sig(2441);
CN_in_sig(3579)	<=	VN_out_sig(2442);
CN_in_sig(4347)	<=	VN_out_sig(2443);
CN_in_sig(987)	<=	VN_out_sig(2444);
CN_in_sig(1947)	<=	VN_out_sig(2445);
CN_in_sig(3587)	<=	VN_out_sig(2446);
CN_in_sig(4355)	<=	VN_out_sig(2447);
CN_in_sig(995)	<=	VN_out_sig(2448);
CN_in_sig(1955)	<=	VN_out_sig(2449);
CN_in_sig(3595)	<=	VN_out_sig(2450);
CN_in_sig(4363)	<=	VN_out_sig(2451);
CN_in_sig(1003)	<=	VN_out_sig(2452);
CN_in_sig(1963)	<=	VN_out_sig(2453);
CN_in_sig(3603)	<=	VN_out_sig(2454);
CN_in_sig(4371)	<=	VN_out_sig(2455);
CN_in_sig(1011)	<=	VN_out_sig(2456);
CN_in_sig(1971)	<=	VN_out_sig(2457);
CN_in_sig(3611)	<=	VN_out_sig(2458);
CN_in_sig(4379)	<=	VN_out_sig(2459);
CN_in_sig(1019)	<=	VN_out_sig(2460);
CN_in_sig(1979)	<=	VN_out_sig(2461);
CN_in_sig(3619)	<=	VN_out_sig(2462);
CN_in_sig(4387)	<=	VN_out_sig(2463);
CN_in_sig(1027)	<=	VN_out_sig(2464);
CN_in_sig(1987)	<=	VN_out_sig(2465);
CN_in_sig(3627)	<=	VN_out_sig(2466);
CN_in_sig(4395)	<=	VN_out_sig(2467);
CN_in_sig(1035)	<=	VN_out_sig(2468);
CN_in_sig(1995)	<=	VN_out_sig(2469);
CN_in_sig(3635)	<=	VN_out_sig(2470);
CN_in_sig(4403)	<=	VN_out_sig(2471);
CN_in_sig(1043)	<=	VN_out_sig(2472);
CN_in_sig(2003)	<=	VN_out_sig(2473);
CN_in_sig(3643)	<=	VN_out_sig(2474);
CN_in_sig(4411)	<=	VN_out_sig(2475);
CN_in_sig(1051)	<=	VN_out_sig(2476);
CN_in_sig(2011)	<=	VN_out_sig(2477);
CN_in_sig(3651)	<=	VN_out_sig(2478);
CN_in_sig(4419)	<=	VN_out_sig(2479);
CN_in_sig(1059)	<=	VN_out_sig(2480);
CN_in_sig(2019)	<=	VN_out_sig(2481);
CN_in_sig(3659)	<=	VN_out_sig(2482);
CN_in_sig(4427)	<=	VN_out_sig(2483);
CN_in_sig(1067)	<=	VN_out_sig(2484);
CN_in_sig(2027)	<=	VN_out_sig(2485);
CN_in_sig(3667)	<=	VN_out_sig(2486);
CN_in_sig(4435)	<=	VN_out_sig(2487);
CN_in_sig(1075)	<=	VN_out_sig(2488);
CN_in_sig(2035)	<=	VN_out_sig(2489);
CN_in_sig(3675)	<=	VN_out_sig(2490);
CN_in_sig(4443)	<=	VN_out_sig(2491);
CN_in_sig(1083)	<=	VN_out_sig(2492);
CN_in_sig(2043)	<=	VN_out_sig(2493);
CN_in_sig(3683)	<=	VN_out_sig(2494);
CN_in_sig(4451)	<=	VN_out_sig(2495);
CN_in_sig(1091)	<=	VN_out_sig(2496);
CN_in_sig(2051)	<=	VN_out_sig(2497);
CN_in_sig(3691)	<=	VN_out_sig(2498);
CN_in_sig(4459)	<=	VN_out_sig(2499);
CN_in_sig(1099)	<=	VN_out_sig(2500);
CN_in_sig(2059)	<=	VN_out_sig(2501);
CN_in_sig(3699)	<=	VN_out_sig(2502);
CN_in_sig(4467)	<=	VN_out_sig(2503);
CN_in_sig(1107)	<=	VN_out_sig(2504);
CN_in_sig(2067)	<=	VN_out_sig(2505);
CN_in_sig(3707)	<=	VN_out_sig(2506);
CN_in_sig(4475)	<=	VN_out_sig(2507);
CN_in_sig(1115)	<=	VN_out_sig(2508);
CN_in_sig(2075)	<=	VN_out_sig(2509);
CN_in_sig(3715)	<=	VN_out_sig(2510);
CN_in_sig(4483)	<=	VN_out_sig(2511);
CN_in_sig(1123)	<=	VN_out_sig(2512);
CN_in_sig(2083)	<=	VN_out_sig(2513);
CN_in_sig(3723)	<=	VN_out_sig(2514);
CN_in_sig(4491)	<=	VN_out_sig(2515);
CN_in_sig(1131)	<=	VN_out_sig(2516);
CN_in_sig(2091)	<=	VN_out_sig(2517);
CN_in_sig(3731)	<=	VN_out_sig(2518);
CN_in_sig(4499)	<=	VN_out_sig(2519);
CN_in_sig(1139)	<=	VN_out_sig(2520);
CN_in_sig(2099)	<=	VN_out_sig(2521);
CN_in_sig(3739)	<=	VN_out_sig(2522);
CN_in_sig(4507)	<=	VN_out_sig(2523);
CN_in_sig(1147)	<=	VN_out_sig(2524);
CN_in_sig(2107)	<=	VN_out_sig(2525);
CN_in_sig(3747)	<=	VN_out_sig(2526);
CN_in_sig(4515)	<=	VN_out_sig(2527);
CN_in_sig(1155)	<=	VN_out_sig(2528);
CN_in_sig(2115)	<=	VN_out_sig(2529);
CN_in_sig(3755)	<=	VN_out_sig(2530);
CN_in_sig(4523)	<=	VN_out_sig(2531);
CN_in_sig(1163)	<=	VN_out_sig(2532);
CN_in_sig(2123)	<=	VN_out_sig(2533);
CN_in_sig(3763)	<=	VN_out_sig(2534);
CN_in_sig(4531)	<=	VN_out_sig(2535);
CN_in_sig(1171)	<=	VN_out_sig(2536);
CN_in_sig(2131)	<=	VN_out_sig(2537);
CN_in_sig(3771)	<=	VN_out_sig(2538);
CN_in_sig(4539)	<=	VN_out_sig(2539);
CN_in_sig(1179)	<=	VN_out_sig(2540);
CN_in_sig(2139)	<=	VN_out_sig(2541);
CN_in_sig(3779)	<=	VN_out_sig(2542);
CN_in_sig(4547)	<=	VN_out_sig(2543);
CN_in_sig(1187)	<=	VN_out_sig(2544);
CN_in_sig(2147)	<=	VN_out_sig(2545);
CN_in_sig(3787)	<=	VN_out_sig(2546);
CN_in_sig(4555)	<=	VN_out_sig(2547);
CN_in_sig(1195)	<=	VN_out_sig(2548);
CN_in_sig(2155)	<=	VN_out_sig(2549);
CN_in_sig(3795)	<=	VN_out_sig(2550);
CN_in_sig(4563)	<=	VN_out_sig(2551);
CN_in_sig(1203)	<=	VN_out_sig(2552);
CN_in_sig(1731)	<=	VN_out_sig(2553);
CN_in_sig(3803)	<=	VN_out_sig(2554);
CN_in_sig(4571)	<=	VN_out_sig(2555);
CN_in_sig(1211)	<=	VN_out_sig(2556);
CN_in_sig(1739)	<=	VN_out_sig(2557);
CN_in_sig(3811)	<=	VN_out_sig(2558);
CN_in_sig(4579)	<=	VN_out_sig(2559);
CN_in_sig(1219)	<=	VN_out_sig(2560);
CN_in_sig(1747)	<=	VN_out_sig(2561);
CN_in_sig(3819)	<=	VN_out_sig(2562);
CN_in_sig(4587)	<=	VN_out_sig(2563);
CN_in_sig(1227)	<=	VN_out_sig(2564);
CN_in_sig(1755)	<=	VN_out_sig(2565);
CN_in_sig(3827)	<=	VN_out_sig(2566);
CN_in_sig(4595)	<=	VN_out_sig(2567);
CN_in_sig(1235)	<=	VN_out_sig(2568);
CN_in_sig(1763)	<=	VN_out_sig(2569);
CN_in_sig(3835)	<=	VN_out_sig(2570);
CN_in_sig(4603)	<=	VN_out_sig(2571);
CN_in_sig(1243)	<=	VN_out_sig(2572);
CN_in_sig(1771)	<=	VN_out_sig(2573);
CN_in_sig(3843)	<=	VN_out_sig(2574);
CN_in_sig(4611)	<=	VN_out_sig(2575);
CN_in_sig(1251)	<=	VN_out_sig(2576);
CN_in_sig(1779)	<=	VN_out_sig(2577);
CN_in_sig(3851)	<=	VN_out_sig(2578);
CN_in_sig(4619)	<=	VN_out_sig(2579);
CN_in_sig(1259)	<=	VN_out_sig(2580);
CN_in_sig(1787)	<=	VN_out_sig(2581);
CN_in_sig(3859)	<=	VN_out_sig(2582);
CN_in_sig(4627)	<=	VN_out_sig(2583);
CN_in_sig(1267)	<=	VN_out_sig(2584);
CN_in_sig(1795)	<=	VN_out_sig(2585);
CN_in_sig(3867)	<=	VN_out_sig(2586);
CN_in_sig(4635)	<=	VN_out_sig(2587);
CN_in_sig(1275)	<=	VN_out_sig(2588);
CN_in_sig(1803)	<=	VN_out_sig(2589);
CN_in_sig(3875)	<=	VN_out_sig(2590);
CN_in_sig(4643)	<=	VN_out_sig(2591);
CN_in_sig(900)	<=	VN_out_sig(2592);
CN_in_sig(2580)	<=	VN_out_sig(2593);
CN_in_sig(3004)	<=	VN_out_sig(2594);
CN_in_sig(4420)	<=	VN_out_sig(2595);
CN_in_sig(908)	<=	VN_out_sig(2596);
CN_in_sig(2588)	<=	VN_out_sig(2597);
CN_in_sig(3012)	<=	VN_out_sig(2598);
CN_in_sig(4428)	<=	VN_out_sig(2599);
CN_in_sig(916)	<=	VN_out_sig(2600);
CN_in_sig(2164)	<=	VN_out_sig(2601);
CN_in_sig(3020)	<=	VN_out_sig(2602);
CN_in_sig(4436)	<=	VN_out_sig(2603);
CN_in_sig(924)	<=	VN_out_sig(2604);
CN_in_sig(2172)	<=	VN_out_sig(2605);
CN_in_sig(2596)	<=	VN_out_sig(2606);
CN_in_sig(4444)	<=	VN_out_sig(2607);
CN_in_sig(932)	<=	VN_out_sig(2608);
CN_in_sig(2180)	<=	VN_out_sig(2609);
CN_in_sig(2604)	<=	VN_out_sig(2610);
CN_in_sig(4452)	<=	VN_out_sig(2611);
CN_in_sig(940)	<=	VN_out_sig(2612);
CN_in_sig(2188)	<=	VN_out_sig(2613);
CN_in_sig(2612)	<=	VN_out_sig(2614);
CN_in_sig(4460)	<=	VN_out_sig(2615);
CN_in_sig(948)	<=	VN_out_sig(2616);
CN_in_sig(2196)	<=	VN_out_sig(2617);
CN_in_sig(2620)	<=	VN_out_sig(2618);
CN_in_sig(4468)	<=	VN_out_sig(2619);
CN_in_sig(956)	<=	VN_out_sig(2620);
CN_in_sig(2204)	<=	VN_out_sig(2621);
CN_in_sig(2628)	<=	VN_out_sig(2622);
CN_in_sig(4476)	<=	VN_out_sig(2623);
CN_in_sig(964)	<=	VN_out_sig(2624);
CN_in_sig(2212)	<=	VN_out_sig(2625);
CN_in_sig(2636)	<=	VN_out_sig(2626);
CN_in_sig(4484)	<=	VN_out_sig(2627);
CN_in_sig(972)	<=	VN_out_sig(2628);
CN_in_sig(2220)	<=	VN_out_sig(2629);
CN_in_sig(2644)	<=	VN_out_sig(2630);
CN_in_sig(4492)	<=	VN_out_sig(2631);
CN_in_sig(980)	<=	VN_out_sig(2632);
CN_in_sig(2228)	<=	VN_out_sig(2633);
CN_in_sig(2652)	<=	VN_out_sig(2634);
CN_in_sig(4500)	<=	VN_out_sig(2635);
CN_in_sig(988)	<=	VN_out_sig(2636);
CN_in_sig(2236)	<=	VN_out_sig(2637);
CN_in_sig(2660)	<=	VN_out_sig(2638);
CN_in_sig(4508)	<=	VN_out_sig(2639);
CN_in_sig(996)	<=	VN_out_sig(2640);
CN_in_sig(2244)	<=	VN_out_sig(2641);
CN_in_sig(2668)	<=	VN_out_sig(2642);
CN_in_sig(4516)	<=	VN_out_sig(2643);
CN_in_sig(1004)	<=	VN_out_sig(2644);
CN_in_sig(2252)	<=	VN_out_sig(2645);
CN_in_sig(2676)	<=	VN_out_sig(2646);
CN_in_sig(4524)	<=	VN_out_sig(2647);
CN_in_sig(1012)	<=	VN_out_sig(2648);
CN_in_sig(2260)	<=	VN_out_sig(2649);
CN_in_sig(2684)	<=	VN_out_sig(2650);
CN_in_sig(4532)	<=	VN_out_sig(2651);
CN_in_sig(1020)	<=	VN_out_sig(2652);
CN_in_sig(2268)	<=	VN_out_sig(2653);
CN_in_sig(2692)	<=	VN_out_sig(2654);
CN_in_sig(4540)	<=	VN_out_sig(2655);
CN_in_sig(1028)	<=	VN_out_sig(2656);
CN_in_sig(2276)	<=	VN_out_sig(2657);
CN_in_sig(2700)	<=	VN_out_sig(2658);
CN_in_sig(4548)	<=	VN_out_sig(2659);
CN_in_sig(1036)	<=	VN_out_sig(2660);
CN_in_sig(2284)	<=	VN_out_sig(2661);
CN_in_sig(2708)	<=	VN_out_sig(2662);
CN_in_sig(4556)	<=	VN_out_sig(2663);
CN_in_sig(1044)	<=	VN_out_sig(2664);
CN_in_sig(2292)	<=	VN_out_sig(2665);
CN_in_sig(2716)	<=	VN_out_sig(2666);
CN_in_sig(4564)	<=	VN_out_sig(2667);
CN_in_sig(1052)	<=	VN_out_sig(2668);
CN_in_sig(2300)	<=	VN_out_sig(2669);
CN_in_sig(2724)	<=	VN_out_sig(2670);
CN_in_sig(4572)	<=	VN_out_sig(2671);
CN_in_sig(1060)	<=	VN_out_sig(2672);
CN_in_sig(2308)	<=	VN_out_sig(2673);
CN_in_sig(2732)	<=	VN_out_sig(2674);
CN_in_sig(4580)	<=	VN_out_sig(2675);
CN_in_sig(1068)	<=	VN_out_sig(2676);
CN_in_sig(2316)	<=	VN_out_sig(2677);
CN_in_sig(2740)	<=	VN_out_sig(2678);
CN_in_sig(4588)	<=	VN_out_sig(2679);
CN_in_sig(1076)	<=	VN_out_sig(2680);
CN_in_sig(2324)	<=	VN_out_sig(2681);
CN_in_sig(2748)	<=	VN_out_sig(2682);
CN_in_sig(4596)	<=	VN_out_sig(2683);
CN_in_sig(1084)	<=	VN_out_sig(2684);
CN_in_sig(2332)	<=	VN_out_sig(2685);
CN_in_sig(2756)	<=	VN_out_sig(2686);
CN_in_sig(4604)	<=	VN_out_sig(2687);
CN_in_sig(1092)	<=	VN_out_sig(2688);
CN_in_sig(2340)	<=	VN_out_sig(2689);
CN_in_sig(2764)	<=	VN_out_sig(2690);
CN_in_sig(4612)	<=	VN_out_sig(2691);
CN_in_sig(1100)	<=	VN_out_sig(2692);
CN_in_sig(2348)	<=	VN_out_sig(2693);
CN_in_sig(2772)	<=	VN_out_sig(2694);
CN_in_sig(4620)	<=	VN_out_sig(2695);
CN_in_sig(1108)	<=	VN_out_sig(2696);
CN_in_sig(2356)	<=	VN_out_sig(2697);
CN_in_sig(2780)	<=	VN_out_sig(2698);
CN_in_sig(4628)	<=	VN_out_sig(2699);
CN_in_sig(1116)	<=	VN_out_sig(2700);
CN_in_sig(2364)	<=	VN_out_sig(2701);
CN_in_sig(2788)	<=	VN_out_sig(2702);
CN_in_sig(4636)	<=	VN_out_sig(2703);
CN_in_sig(1124)	<=	VN_out_sig(2704);
CN_in_sig(2372)	<=	VN_out_sig(2705);
CN_in_sig(2796)	<=	VN_out_sig(2706);
CN_in_sig(4644)	<=	VN_out_sig(2707);
CN_in_sig(1132)	<=	VN_out_sig(2708);
CN_in_sig(2380)	<=	VN_out_sig(2709);
CN_in_sig(2804)	<=	VN_out_sig(2710);
CN_in_sig(4652)	<=	VN_out_sig(2711);
CN_in_sig(1140)	<=	VN_out_sig(2712);
CN_in_sig(2388)	<=	VN_out_sig(2713);
CN_in_sig(2812)	<=	VN_out_sig(2714);
CN_in_sig(4660)	<=	VN_out_sig(2715);
CN_in_sig(1148)	<=	VN_out_sig(2716);
CN_in_sig(2396)	<=	VN_out_sig(2717);
CN_in_sig(2820)	<=	VN_out_sig(2718);
CN_in_sig(4668)	<=	VN_out_sig(2719);
CN_in_sig(1156)	<=	VN_out_sig(2720);
CN_in_sig(2404)	<=	VN_out_sig(2721);
CN_in_sig(2828)	<=	VN_out_sig(2722);
CN_in_sig(4676)	<=	VN_out_sig(2723);
CN_in_sig(1164)	<=	VN_out_sig(2724);
CN_in_sig(2412)	<=	VN_out_sig(2725);
CN_in_sig(2836)	<=	VN_out_sig(2726);
CN_in_sig(4684)	<=	VN_out_sig(2727);
CN_in_sig(1172)	<=	VN_out_sig(2728);
CN_in_sig(2420)	<=	VN_out_sig(2729);
CN_in_sig(2844)	<=	VN_out_sig(2730);
CN_in_sig(4692)	<=	VN_out_sig(2731);
CN_in_sig(1180)	<=	VN_out_sig(2732);
CN_in_sig(2428)	<=	VN_out_sig(2733);
CN_in_sig(2852)	<=	VN_out_sig(2734);
CN_in_sig(4700)	<=	VN_out_sig(2735);
CN_in_sig(1188)	<=	VN_out_sig(2736);
CN_in_sig(2436)	<=	VN_out_sig(2737);
CN_in_sig(2860)	<=	VN_out_sig(2738);
CN_in_sig(4708)	<=	VN_out_sig(2739);
CN_in_sig(1196)	<=	VN_out_sig(2740);
CN_in_sig(2444)	<=	VN_out_sig(2741);
CN_in_sig(2868)	<=	VN_out_sig(2742);
CN_in_sig(4716)	<=	VN_out_sig(2743);
CN_in_sig(1204)	<=	VN_out_sig(2744);
CN_in_sig(2452)	<=	VN_out_sig(2745);
CN_in_sig(2876)	<=	VN_out_sig(2746);
CN_in_sig(4724)	<=	VN_out_sig(2747);
CN_in_sig(1212)	<=	VN_out_sig(2748);
CN_in_sig(2460)	<=	VN_out_sig(2749);
CN_in_sig(2884)	<=	VN_out_sig(2750);
CN_in_sig(4732)	<=	VN_out_sig(2751);
CN_in_sig(1220)	<=	VN_out_sig(2752);
CN_in_sig(2468)	<=	VN_out_sig(2753);
CN_in_sig(2892)	<=	VN_out_sig(2754);
CN_in_sig(4740)	<=	VN_out_sig(2755);
CN_in_sig(1228)	<=	VN_out_sig(2756);
CN_in_sig(2476)	<=	VN_out_sig(2757);
CN_in_sig(2900)	<=	VN_out_sig(2758);
CN_in_sig(4748)	<=	VN_out_sig(2759);
CN_in_sig(1236)	<=	VN_out_sig(2760);
CN_in_sig(2484)	<=	VN_out_sig(2761);
CN_in_sig(2908)	<=	VN_out_sig(2762);
CN_in_sig(4324)	<=	VN_out_sig(2763);
CN_in_sig(1244)	<=	VN_out_sig(2764);
CN_in_sig(2492)	<=	VN_out_sig(2765);
CN_in_sig(2916)	<=	VN_out_sig(2766);
CN_in_sig(4332)	<=	VN_out_sig(2767);
CN_in_sig(1252)	<=	VN_out_sig(2768);
CN_in_sig(2500)	<=	VN_out_sig(2769);
CN_in_sig(2924)	<=	VN_out_sig(2770);
CN_in_sig(4340)	<=	VN_out_sig(2771);
CN_in_sig(1260)	<=	VN_out_sig(2772);
CN_in_sig(2508)	<=	VN_out_sig(2773);
CN_in_sig(2932)	<=	VN_out_sig(2774);
CN_in_sig(4348)	<=	VN_out_sig(2775);
CN_in_sig(1268)	<=	VN_out_sig(2776);
CN_in_sig(2516)	<=	VN_out_sig(2777);
CN_in_sig(2940)	<=	VN_out_sig(2778);
CN_in_sig(4356)	<=	VN_out_sig(2779);
CN_in_sig(1276)	<=	VN_out_sig(2780);
CN_in_sig(2524)	<=	VN_out_sig(2781);
CN_in_sig(2948)	<=	VN_out_sig(2782);
CN_in_sig(4364)	<=	VN_out_sig(2783);
CN_in_sig(1284)	<=	VN_out_sig(2784);
CN_in_sig(2532)	<=	VN_out_sig(2785);
CN_in_sig(2956)	<=	VN_out_sig(2786);
CN_in_sig(4372)	<=	VN_out_sig(2787);
CN_in_sig(1292)	<=	VN_out_sig(2788);
CN_in_sig(2540)	<=	VN_out_sig(2789);
CN_in_sig(2964)	<=	VN_out_sig(2790);
CN_in_sig(4380)	<=	VN_out_sig(2791);
CN_in_sig(868)	<=	VN_out_sig(2792);
CN_in_sig(2548)	<=	VN_out_sig(2793);
CN_in_sig(2972)	<=	VN_out_sig(2794);
CN_in_sig(4388)	<=	VN_out_sig(2795);
CN_in_sig(876)	<=	VN_out_sig(2796);
CN_in_sig(2556)	<=	VN_out_sig(2797);
CN_in_sig(2980)	<=	VN_out_sig(2798);
CN_in_sig(4396)	<=	VN_out_sig(2799);
CN_in_sig(884)	<=	VN_out_sig(2800);
CN_in_sig(2564)	<=	VN_out_sig(2801);
CN_in_sig(2988)	<=	VN_out_sig(2802);
CN_in_sig(4404)	<=	VN_out_sig(2803);
CN_in_sig(892)	<=	VN_out_sig(2804);
CN_in_sig(2572)	<=	VN_out_sig(2805);
CN_in_sig(2996)	<=	VN_out_sig(2806);
CN_in_sig(4412)	<=	VN_out_sig(2807);
CN_in_sig(84)	<=	VN_out_sig(2808);
CN_in_sig(1628)	<=	VN_out_sig(2809);
CN_in_sig(3740)	<=	VN_out_sig(2810);
CN_in_sig(4820)	<=	VN_out_sig(2811);
CN_in_sig(92)	<=	VN_out_sig(2812);
CN_in_sig(1636)	<=	VN_out_sig(2813);
CN_in_sig(3748)	<=	VN_out_sig(2814);
CN_in_sig(4828)	<=	VN_out_sig(2815);
CN_in_sig(100)	<=	VN_out_sig(2816);
CN_in_sig(1644)	<=	VN_out_sig(2817);
CN_in_sig(3756)	<=	VN_out_sig(2818);
CN_in_sig(4836)	<=	VN_out_sig(2819);
CN_in_sig(108)	<=	VN_out_sig(2820);
CN_in_sig(1652)	<=	VN_out_sig(2821);
CN_in_sig(3764)	<=	VN_out_sig(2822);
CN_in_sig(4844)	<=	VN_out_sig(2823);
CN_in_sig(116)	<=	VN_out_sig(2824);
CN_in_sig(1660)	<=	VN_out_sig(2825);
CN_in_sig(3772)	<=	VN_out_sig(2826);
CN_in_sig(4852)	<=	VN_out_sig(2827);
CN_in_sig(124)	<=	VN_out_sig(2828);
CN_in_sig(1668)	<=	VN_out_sig(2829);
CN_in_sig(3780)	<=	VN_out_sig(2830);
CN_in_sig(4860)	<=	VN_out_sig(2831);
CN_in_sig(132)	<=	VN_out_sig(2832);
CN_in_sig(1676)	<=	VN_out_sig(2833);
CN_in_sig(3788)	<=	VN_out_sig(2834);
CN_in_sig(4868)	<=	VN_out_sig(2835);
CN_in_sig(140)	<=	VN_out_sig(2836);
CN_in_sig(1684)	<=	VN_out_sig(2837);
CN_in_sig(3796)	<=	VN_out_sig(2838);
CN_in_sig(4876)	<=	VN_out_sig(2839);
CN_in_sig(148)	<=	VN_out_sig(2840);
CN_in_sig(1692)	<=	VN_out_sig(2841);
CN_in_sig(3804)	<=	VN_out_sig(2842);
CN_in_sig(4884)	<=	VN_out_sig(2843);
CN_in_sig(156)	<=	VN_out_sig(2844);
CN_in_sig(1700)	<=	VN_out_sig(2845);
CN_in_sig(3812)	<=	VN_out_sig(2846);
CN_in_sig(4892)	<=	VN_out_sig(2847);
CN_in_sig(164)	<=	VN_out_sig(2848);
CN_in_sig(1708)	<=	VN_out_sig(2849);
CN_in_sig(3820)	<=	VN_out_sig(2850);
CN_in_sig(4900)	<=	VN_out_sig(2851);
CN_in_sig(172)	<=	VN_out_sig(2852);
CN_in_sig(1716)	<=	VN_out_sig(2853);
CN_in_sig(3828)	<=	VN_out_sig(2854);
CN_in_sig(4908)	<=	VN_out_sig(2855);
CN_in_sig(180)	<=	VN_out_sig(2856);
CN_in_sig(1724)	<=	VN_out_sig(2857);
CN_in_sig(3836)	<=	VN_out_sig(2858);
CN_in_sig(4916)	<=	VN_out_sig(2859);
CN_in_sig(188)	<=	VN_out_sig(2860);
CN_in_sig(1300)	<=	VN_out_sig(2861);
CN_in_sig(3844)	<=	VN_out_sig(2862);
CN_in_sig(4924)	<=	VN_out_sig(2863);
CN_in_sig(196)	<=	VN_out_sig(2864);
CN_in_sig(1308)	<=	VN_out_sig(2865);
CN_in_sig(3852)	<=	VN_out_sig(2866);
CN_in_sig(4932)	<=	VN_out_sig(2867);
CN_in_sig(204)	<=	VN_out_sig(2868);
CN_in_sig(1316)	<=	VN_out_sig(2869);
CN_in_sig(3860)	<=	VN_out_sig(2870);
CN_in_sig(4940)	<=	VN_out_sig(2871);
CN_in_sig(212)	<=	VN_out_sig(2872);
CN_in_sig(1324)	<=	VN_out_sig(2873);
CN_in_sig(3868)	<=	VN_out_sig(2874);
CN_in_sig(4948)	<=	VN_out_sig(2875);
CN_in_sig(220)	<=	VN_out_sig(2876);
CN_in_sig(1332)	<=	VN_out_sig(2877);
CN_in_sig(3876)	<=	VN_out_sig(2878);
CN_in_sig(4956)	<=	VN_out_sig(2879);
CN_in_sig(228)	<=	VN_out_sig(2880);
CN_in_sig(1340)	<=	VN_out_sig(2881);
CN_in_sig(3884)	<=	VN_out_sig(2882);
CN_in_sig(4964)	<=	VN_out_sig(2883);
CN_in_sig(236)	<=	VN_out_sig(2884);
CN_in_sig(1348)	<=	VN_out_sig(2885);
CN_in_sig(3460)	<=	VN_out_sig(2886);
CN_in_sig(4972)	<=	VN_out_sig(2887);
CN_in_sig(244)	<=	VN_out_sig(2888);
CN_in_sig(1356)	<=	VN_out_sig(2889);
CN_in_sig(3468)	<=	VN_out_sig(2890);
CN_in_sig(4980)	<=	VN_out_sig(2891);
CN_in_sig(252)	<=	VN_out_sig(2892);
CN_in_sig(1364)	<=	VN_out_sig(2893);
CN_in_sig(3476)	<=	VN_out_sig(2894);
CN_in_sig(4988)	<=	VN_out_sig(2895);
CN_in_sig(260)	<=	VN_out_sig(2896);
CN_in_sig(1372)	<=	VN_out_sig(2897);
CN_in_sig(3484)	<=	VN_out_sig(2898);
CN_in_sig(4996)	<=	VN_out_sig(2899);
CN_in_sig(268)	<=	VN_out_sig(2900);
CN_in_sig(1380)	<=	VN_out_sig(2901);
CN_in_sig(3492)	<=	VN_out_sig(2902);
CN_in_sig(5004)	<=	VN_out_sig(2903);
CN_in_sig(276)	<=	VN_out_sig(2904);
CN_in_sig(1388)	<=	VN_out_sig(2905);
CN_in_sig(3500)	<=	VN_out_sig(2906);
CN_in_sig(5012)	<=	VN_out_sig(2907);
CN_in_sig(284)	<=	VN_out_sig(2908);
CN_in_sig(1396)	<=	VN_out_sig(2909);
CN_in_sig(3508)	<=	VN_out_sig(2910);
CN_in_sig(5020)	<=	VN_out_sig(2911);
CN_in_sig(292)	<=	VN_out_sig(2912);
CN_in_sig(1404)	<=	VN_out_sig(2913);
CN_in_sig(3516)	<=	VN_out_sig(2914);
CN_in_sig(5028)	<=	VN_out_sig(2915);
CN_in_sig(300)	<=	VN_out_sig(2916);
CN_in_sig(1412)	<=	VN_out_sig(2917);
CN_in_sig(3524)	<=	VN_out_sig(2918);
CN_in_sig(5036)	<=	VN_out_sig(2919);
CN_in_sig(308)	<=	VN_out_sig(2920);
CN_in_sig(1420)	<=	VN_out_sig(2921);
CN_in_sig(3532)	<=	VN_out_sig(2922);
CN_in_sig(5044)	<=	VN_out_sig(2923);
CN_in_sig(316)	<=	VN_out_sig(2924);
CN_in_sig(1428)	<=	VN_out_sig(2925);
CN_in_sig(3540)	<=	VN_out_sig(2926);
CN_in_sig(5052)	<=	VN_out_sig(2927);
CN_in_sig(324)	<=	VN_out_sig(2928);
CN_in_sig(1436)	<=	VN_out_sig(2929);
CN_in_sig(3548)	<=	VN_out_sig(2930);
CN_in_sig(5060)	<=	VN_out_sig(2931);
CN_in_sig(332)	<=	VN_out_sig(2932);
CN_in_sig(1444)	<=	VN_out_sig(2933);
CN_in_sig(3556)	<=	VN_out_sig(2934);
CN_in_sig(5068)	<=	VN_out_sig(2935);
CN_in_sig(340)	<=	VN_out_sig(2936);
CN_in_sig(1452)	<=	VN_out_sig(2937);
CN_in_sig(3564)	<=	VN_out_sig(2938);
CN_in_sig(5076)	<=	VN_out_sig(2939);
CN_in_sig(348)	<=	VN_out_sig(2940);
CN_in_sig(1460)	<=	VN_out_sig(2941);
CN_in_sig(3572)	<=	VN_out_sig(2942);
CN_in_sig(5084)	<=	VN_out_sig(2943);
CN_in_sig(356)	<=	VN_out_sig(2944);
CN_in_sig(1468)	<=	VN_out_sig(2945);
CN_in_sig(3580)	<=	VN_out_sig(2946);
CN_in_sig(5092)	<=	VN_out_sig(2947);
CN_in_sig(364)	<=	VN_out_sig(2948);
CN_in_sig(1476)	<=	VN_out_sig(2949);
CN_in_sig(3588)	<=	VN_out_sig(2950);
CN_in_sig(5100)	<=	VN_out_sig(2951);
CN_in_sig(372)	<=	VN_out_sig(2952);
CN_in_sig(1484)	<=	VN_out_sig(2953);
CN_in_sig(3596)	<=	VN_out_sig(2954);
CN_in_sig(5108)	<=	VN_out_sig(2955);
CN_in_sig(380)	<=	VN_out_sig(2956);
CN_in_sig(1492)	<=	VN_out_sig(2957);
CN_in_sig(3604)	<=	VN_out_sig(2958);
CN_in_sig(5116)	<=	VN_out_sig(2959);
CN_in_sig(388)	<=	VN_out_sig(2960);
CN_in_sig(1500)	<=	VN_out_sig(2961);
CN_in_sig(3612)	<=	VN_out_sig(2962);
CN_in_sig(5124)	<=	VN_out_sig(2963);
CN_in_sig(396)	<=	VN_out_sig(2964);
CN_in_sig(1508)	<=	VN_out_sig(2965);
CN_in_sig(3620)	<=	VN_out_sig(2966);
CN_in_sig(5132)	<=	VN_out_sig(2967);
CN_in_sig(404)	<=	VN_out_sig(2968);
CN_in_sig(1516)	<=	VN_out_sig(2969);
CN_in_sig(3628)	<=	VN_out_sig(2970);
CN_in_sig(5140)	<=	VN_out_sig(2971);
CN_in_sig(412)	<=	VN_out_sig(2972);
CN_in_sig(1524)	<=	VN_out_sig(2973);
CN_in_sig(3636)	<=	VN_out_sig(2974);
CN_in_sig(5148)	<=	VN_out_sig(2975);
CN_in_sig(420)	<=	VN_out_sig(2976);
CN_in_sig(1532)	<=	VN_out_sig(2977);
CN_in_sig(3644)	<=	VN_out_sig(2978);
CN_in_sig(5156)	<=	VN_out_sig(2979);
CN_in_sig(428)	<=	VN_out_sig(2980);
CN_in_sig(1540)	<=	VN_out_sig(2981);
CN_in_sig(3652)	<=	VN_out_sig(2982);
CN_in_sig(5164)	<=	VN_out_sig(2983);
CN_in_sig(4)	<=	VN_out_sig(2984);
CN_in_sig(1548)	<=	VN_out_sig(2985);
CN_in_sig(3660)	<=	VN_out_sig(2986);
CN_in_sig(5172)	<=	VN_out_sig(2987);
CN_in_sig(12)	<=	VN_out_sig(2988);
CN_in_sig(1556)	<=	VN_out_sig(2989);
CN_in_sig(3668)	<=	VN_out_sig(2990);
CN_in_sig(5180)	<=	VN_out_sig(2991);
CN_in_sig(20)	<=	VN_out_sig(2992);
CN_in_sig(1564)	<=	VN_out_sig(2993);
CN_in_sig(3676)	<=	VN_out_sig(2994);
CN_in_sig(4756)	<=	VN_out_sig(2995);
CN_in_sig(28)	<=	VN_out_sig(2996);
CN_in_sig(1572)	<=	VN_out_sig(2997);
CN_in_sig(3684)	<=	VN_out_sig(2998);
CN_in_sig(4764)	<=	VN_out_sig(2999);
CN_in_sig(36)	<=	VN_out_sig(3000);
CN_in_sig(1580)	<=	VN_out_sig(3001);
CN_in_sig(3692)	<=	VN_out_sig(3002);
CN_in_sig(4772)	<=	VN_out_sig(3003);
CN_in_sig(44)	<=	VN_out_sig(3004);
CN_in_sig(1588)	<=	VN_out_sig(3005);
CN_in_sig(3700)	<=	VN_out_sig(3006);
CN_in_sig(4780)	<=	VN_out_sig(3007);
CN_in_sig(52)	<=	VN_out_sig(3008);
CN_in_sig(1596)	<=	VN_out_sig(3009);
CN_in_sig(3708)	<=	VN_out_sig(3010);
CN_in_sig(4788)	<=	VN_out_sig(3011);
CN_in_sig(60)	<=	VN_out_sig(3012);
CN_in_sig(1604)	<=	VN_out_sig(3013);
CN_in_sig(3716)	<=	VN_out_sig(3014);
CN_in_sig(4796)	<=	VN_out_sig(3015);
CN_in_sig(68)	<=	VN_out_sig(3016);
CN_in_sig(1612)	<=	VN_out_sig(3017);
CN_in_sig(3724)	<=	VN_out_sig(3018);
CN_in_sig(4804)	<=	VN_out_sig(3019);
CN_in_sig(76)	<=	VN_out_sig(3020);
CN_in_sig(1620)	<=	VN_out_sig(3021);
CN_in_sig(3732)	<=	VN_out_sig(3022);
CN_in_sig(4812)	<=	VN_out_sig(3023);
CN_in_sig(580)	<=	VN_out_sig(3024);
CN_in_sig(2132)	<=	VN_out_sig(3025);
CN_in_sig(3084)	<=	VN_out_sig(3026);
CN_in_sig(4084)	<=	VN_out_sig(3027);
CN_in_sig(588)	<=	VN_out_sig(3028);
CN_in_sig(2140)	<=	VN_out_sig(3029);
CN_in_sig(3092)	<=	VN_out_sig(3030);
CN_in_sig(4092)	<=	VN_out_sig(3031);
CN_in_sig(596)	<=	VN_out_sig(3032);
CN_in_sig(2148)	<=	VN_out_sig(3033);
CN_in_sig(3100)	<=	VN_out_sig(3034);
CN_in_sig(4100)	<=	VN_out_sig(3035);
CN_in_sig(604)	<=	VN_out_sig(3036);
CN_in_sig(2156)	<=	VN_out_sig(3037);
CN_in_sig(3108)	<=	VN_out_sig(3038);
CN_in_sig(4108)	<=	VN_out_sig(3039);
CN_in_sig(612)	<=	VN_out_sig(3040);
CN_in_sig(1732)	<=	VN_out_sig(3041);
CN_in_sig(3116)	<=	VN_out_sig(3042);
CN_in_sig(4116)	<=	VN_out_sig(3043);
CN_in_sig(620)	<=	VN_out_sig(3044);
CN_in_sig(1740)	<=	VN_out_sig(3045);
CN_in_sig(3124)	<=	VN_out_sig(3046);
CN_in_sig(4124)	<=	VN_out_sig(3047);
CN_in_sig(628)	<=	VN_out_sig(3048);
CN_in_sig(1748)	<=	VN_out_sig(3049);
CN_in_sig(3132)	<=	VN_out_sig(3050);
CN_in_sig(4132)	<=	VN_out_sig(3051);
CN_in_sig(636)	<=	VN_out_sig(3052);
CN_in_sig(1756)	<=	VN_out_sig(3053);
CN_in_sig(3140)	<=	VN_out_sig(3054);
CN_in_sig(4140)	<=	VN_out_sig(3055);
CN_in_sig(644)	<=	VN_out_sig(3056);
CN_in_sig(1764)	<=	VN_out_sig(3057);
CN_in_sig(3148)	<=	VN_out_sig(3058);
CN_in_sig(4148)	<=	VN_out_sig(3059);
CN_in_sig(652)	<=	VN_out_sig(3060);
CN_in_sig(1772)	<=	VN_out_sig(3061);
CN_in_sig(3156)	<=	VN_out_sig(3062);
CN_in_sig(4156)	<=	VN_out_sig(3063);
CN_in_sig(660)	<=	VN_out_sig(3064);
CN_in_sig(1780)	<=	VN_out_sig(3065);
CN_in_sig(3164)	<=	VN_out_sig(3066);
CN_in_sig(4164)	<=	VN_out_sig(3067);
CN_in_sig(668)	<=	VN_out_sig(3068);
CN_in_sig(1788)	<=	VN_out_sig(3069);
CN_in_sig(3172)	<=	VN_out_sig(3070);
CN_in_sig(4172)	<=	VN_out_sig(3071);
CN_in_sig(676)	<=	VN_out_sig(3072);
CN_in_sig(1796)	<=	VN_out_sig(3073);
CN_in_sig(3180)	<=	VN_out_sig(3074);
CN_in_sig(4180)	<=	VN_out_sig(3075);
CN_in_sig(684)	<=	VN_out_sig(3076);
CN_in_sig(1804)	<=	VN_out_sig(3077);
CN_in_sig(3188)	<=	VN_out_sig(3078);
CN_in_sig(4188)	<=	VN_out_sig(3079);
CN_in_sig(692)	<=	VN_out_sig(3080);
CN_in_sig(1812)	<=	VN_out_sig(3081);
CN_in_sig(3196)	<=	VN_out_sig(3082);
CN_in_sig(4196)	<=	VN_out_sig(3083);
CN_in_sig(700)	<=	VN_out_sig(3084);
CN_in_sig(1820)	<=	VN_out_sig(3085);
CN_in_sig(3204)	<=	VN_out_sig(3086);
CN_in_sig(4204)	<=	VN_out_sig(3087);
CN_in_sig(708)	<=	VN_out_sig(3088);
CN_in_sig(1828)	<=	VN_out_sig(3089);
CN_in_sig(3212)	<=	VN_out_sig(3090);
CN_in_sig(4212)	<=	VN_out_sig(3091);
CN_in_sig(716)	<=	VN_out_sig(3092);
CN_in_sig(1836)	<=	VN_out_sig(3093);
CN_in_sig(3220)	<=	VN_out_sig(3094);
CN_in_sig(4220)	<=	VN_out_sig(3095);
CN_in_sig(724)	<=	VN_out_sig(3096);
CN_in_sig(1844)	<=	VN_out_sig(3097);
CN_in_sig(3228)	<=	VN_out_sig(3098);
CN_in_sig(4228)	<=	VN_out_sig(3099);
CN_in_sig(732)	<=	VN_out_sig(3100);
CN_in_sig(1852)	<=	VN_out_sig(3101);
CN_in_sig(3236)	<=	VN_out_sig(3102);
CN_in_sig(4236)	<=	VN_out_sig(3103);
CN_in_sig(740)	<=	VN_out_sig(3104);
CN_in_sig(1860)	<=	VN_out_sig(3105);
CN_in_sig(3244)	<=	VN_out_sig(3106);
CN_in_sig(4244)	<=	VN_out_sig(3107);
CN_in_sig(748)	<=	VN_out_sig(3108);
CN_in_sig(1868)	<=	VN_out_sig(3109);
CN_in_sig(3252)	<=	VN_out_sig(3110);
CN_in_sig(4252)	<=	VN_out_sig(3111);
CN_in_sig(756)	<=	VN_out_sig(3112);
CN_in_sig(1876)	<=	VN_out_sig(3113);
CN_in_sig(3260)	<=	VN_out_sig(3114);
CN_in_sig(4260)	<=	VN_out_sig(3115);
CN_in_sig(764)	<=	VN_out_sig(3116);
CN_in_sig(1884)	<=	VN_out_sig(3117);
CN_in_sig(3268)	<=	VN_out_sig(3118);
CN_in_sig(4268)	<=	VN_out_sig(3119);
CN_in_sig(772)	<=	VN_out_sig(3120);
CN_in_sig(1892)	<=	VN_out_sig(3121);
CN_in_sig(3276)	<=	VN_out_sig(3122);
CN_in_sig(4276)	<=	VN_out_sig(3123);
CN_in_sig(780)	<=	VN_out_sig(3124);
CN_in_sig(1900)	<=	VN_out_sig(3125);
CN_in_sig(3284)	<=	VN_out_sig(3126);
CN_in_sig(4284)	<=	VN_out_sig(3127);
CN_in_sig(788)	<=	VN_out_sig(3128);
CN_in_sig(1908)	<=	VN_out_sig(3129);
CN_in_sig(3292)	<=	VN_out_sig(3130);
CN_in_sig(4292)	<=	VN_out_sig(3131);
CN_in_sig(796)	<=	VN_out_sig(3132);
CN_in_sig(1916)	<=	VN_out_sig(3133);
CN_in_sig(3300)	<=	VN_out_sig(3134);
CN_in_sig(4300)	<=	VN_out_sig(3135);
CN_in_sig(804)	<=	VN_out_sig(3136);
CN_in_sig(1924)	<=	VN_out_sig(3137);
CN_in_sig(3308)	<=	VN_out_sig(3138);
CN_in_sig(4308)	<=	VN_out_sig(3139);
CN_in_sig(812)	<=	VN_out_sig(3140);
CN_in_sig(1932)	<=	VN_out_sig(3141);
CN_in_sig(3316)	<=	VN_out_sig(3142);
CN_in_sig(4316)	<=	VN_out_sig(3143);
CN_in_sig(820)	<=	VN_out_sig(3144);
CN_in_sig(1940)	<=	VN_out_sig(3145);
CN_in_sig(3324)	<=	VN_out_sig(3146);
CN_in_sig(3892)	<=	VN_out_sig(3147);
CN_in_sig(828)	<=	VN_out_sig(3148);
CN_in_sig(1948)	<=	VN_out_sig(3149);
CN_in_sig(3332)	<=	VN_out_sig(3150);
CN_in_sig(3900)	<=	VN_out_sig(3151);
CN_in_sig(836)	<=	VN_out_sig(3152);
CN_in_sig(1956)	<=	VN_out_sig(3153);
CN_in_sig(3340)	<=	VN_out_sig(3154);
CN_in_sig(3908)	<=	VN_out_sig(3155);
CN_in_sig(844)	<=	VN_out_sig(3156);
CN_in_sig(1964)	<=	VN_out_sig(3157);
CN_in_sig(3348)	<=	VN_out_sig(3158);
CN_in_sig(3916)	<=	VN_out_sig(3159);
CN_in_sig(852)	<=	VN_out_sig(3160);
CN_in_sig(1972)	<=	VN_out_sig(3161);
CN_in_sig(3356)	<=	VN_out_sig(3162);
CN_in_sig(3924)	<=	VN_out_sig(3163);
CN_in_sig(860)	<=	VN_out_sig(3164);
CN_in_sig(1980)	<=	VN_out_sig(3165);
CN_in_sig(3364)	<=	VN_out_sig(3166);
CN_in_sig(3932)	<=	VN_out_sig(3167);
CN_in_sig(436)	<=	VN_out_sig(3168);
CN_in_sig(1988)	<=	VN_out_sig(3169);
CN_in_sig(3372)	<=	VN_out_sig(3170);
CN_in_sig(3940)	<=	VN_out_sig(3171);
CN_in_sig(444)	<=	VN_out_sig(3172);
CN_in_sig(1996)	<=	VN_out_sig(3173);
CN_in_sig(3380)	<=	VN_out_sig(3174);
CN_in_sig(3948)	<=	VN_out_sig(3175);
CN_in_sig(452)	<=	VN_out_sig(3176);
CN_in_sig(2004)	<=	VN_out_sig(3177);
CN_in_sig(3388)	<=	VN_out_sig(3178);
CN_in_sig(3956)	<=	VN_out_sig(3179);
CN_in_sig(460)	<=	VN_out_sig(3180);
CN_in_sig(2012)	<=	VN_out_sig(3181);
CN_in_sig(3396)	<=	VN_out_sig(3182);
CN_in_sig(3964)	<=	VN_out_sig(3183);
CN_in_sig(468)	<=	VN_out_sig(3184);
CN_in_sig(2020)	<=	VN_out_sig(3185);
CN_in_sig(3404)	<=	VN_out_sig(3186);
CN_in_sig(3972)	<=	VN_out_sig(3187);
CN_in_sig(476)	<=	VN_out_sig(3188);
CN_in_sig(2028)	<=	VN_out_sig(3189);
CN_in_sig(3412)	<=	VN_out_sig(3190);
CN_in_sig(3980)	<=	VN_out_sig(3191);
CN_in_sig(484)	<=	VN_out_sig(3192);
CN_in_sig(2036)	<=	VN_out_sig(3193);
CN_in_sig(3420)	<=	VN_out_sig(3194);
CN_in_sig(3988)	<=	VN_out_sig(3195);
CN_in_sig(492)	<=	VN_out_sig(3196);
CN_in_sig(2044)	<=	VN_out_sig(3197);
CN_in_sig(3428)	<=	VN_out_sig(3198);
CN_in_sig(3996)	<=	VN_out_sig(3199);
CN_in_sig(500)	<=	VN_out_sig(3200);
CN_in_sig(2052)	<=	VN_out_sig(3201);
CN_in_sig(3436)	<=	VN_out_sig(3202);
CN_in_sig(4004)	<=	VN_out_sig(3203);
CN_in_sig(508)	<=	VN_out_sig(3204);
CN_in_sig(2060)	<=	VN_out_sig(3205);
CN_in_sig(3444)	<=	VN_out_sig(3206);
CN_in_sig(4012)	<=	VN_out_sig(3207);
CN_in_sig(516)	<=	VN_out_sig(3208);
CN_in_sig(2068)	<=	VN_out_sig(3209);
CN_in_sig(3452)	<=	VN_out_sig(3210);
CN_in_sig(4020)	<=	VN_out_sig(3211);
CN_in_sig(524)	<=	VN_out_sig(3212);
CN_in_sig(2076)	<=	VN_out_sig(3213);
CN_in_sig(3028)	<=	VN_out_sig(3214);
CN_in_sig(4028)	<=	VN_out_sig(3215);
CN_in_sig(532)	<=	VN_out_sig(3216);
CN_in_sig(2084)	<=	VN_out_sig(3217);
CN_in_sig(3036)	<=	VN_out_sig(3218);
CN_in_sig(4036)	<=	VN_out_sig(3219);
CN_in_sig(540)	<=	VN_out_sig(3220);
CN_in_sig(2092)	<=	VN_out_sig(3221);
CN_in_sig(3044)	<=	VN_out_sig(3222);
CN_in_sig(4044)	<=	VN_out_sig(3223);
CN_in_sig(548)	<=	VN_out_sig(3224);
CN_in_sig(2100)	<=	VN_out_sig(3225);
CN_in_sig(3052)	<=	VN_out_sig(3226);
CN_in_sig(4052)	<=	VN_out_sig(3227);
CN_in_sig(556)	<=	VN_out_sig(3228);
CN_in_sig(2108)	<=	VN_out_sig(3229);
CN_in_sig(3060)	<=	VN_out_sig(3230);
CN_in_sig(4060)	<=	VN_out_sig(3231);
CN_in_sig(564)	<=	VN_out_sig(3232);
CN_in_sig(2116)	<=	VN_out_sig(3233);
CN_in_sig(3068)	<=	VN_out_sig(3234);
CN_in_sig(4068)	<=	VN_out_sig(3235);
CN_in_sig(572)	<=	VN_out_sig(3236);
CN_in_sig(2124)	<=	VN_out_sig(3237);
CN_in_sig(3076)	<=	VN_out_sig(3238);
CN_in_sig(4076)	<=	VN_out_sig(3239);
CN_in_sig(885)	<=	VN_out_sig(3240);
CN_in_sig(2053)	<=	VN_out_sig(3241);
CN_in_sig(2693)	<=	VN_out_sig(3242);
CN_in_sig(4357)	<=	VN_out_sig(3243);
CN_in_sig(893)	<=	VN_out_sig(3244);
CN_in_sig(2061)	<=	VN_out_sig(3245);
CN_in_sig(2701)	<=	VN_out_sig(3246);
CN_in_sig(4365)	<=	VN_out_sig(3247);
CN_in_sig(901)	<=	VN_out_sig(3248);
CN_in_sig(2069)	<=	VN_out_sig(3249);
CN_in_sig(2709)	<=	VN_out_sig(3250);
CN_in_sig(4373)	<=	VN_out_sig(3251);
CN_in_sig(909)	<=	VN_out_sig(3252);
CN_in_sig(2077)	<=	VN_out_sig(3253);
CN_in_sig(2717)	<=	VN_out_sig(3254);
CN_in_sig(4381)	<=	VN_out_sig(3255);
CN_in_sig(917)	<=	VN_out_sig(3256);
CN_in_sig(2085)	<=	VN_out_sig(3257);
CN_in_sig(2725)	<=	VN_out_sig(3258);
CN_in_sig(4389)	<=	VN_out_sig(3259);
CN_in_sig(925)	<=	VN_out_sig(3260);
CN_in_sig(2093)	<=	VN_out_sig(3261);
CN_in_sig(2733)	<=	VN_out_sig(3262);
CN_in_sig(4397)	<=	VN_out_sig(3263);
CN_in_sig(933)	<=	VN_out_sig(3264);
CN_in_sig(2101)	<=	VN_out_sig(3265);
CN_in_sig(2741)	<=	VN_out_sig(3266);
CN_in_sig(4405)	<=	VN_out_sig(3267);
CN_in_sig(941)	<=	VN_out_sig(3268);
CN_in_sig(2109)	<=	VN_out_sig(3269);
CN_in_sig(2749)	<=	VN_out_sig(3270);
CN_in_sig(4413)	<=	VN_out_sig(3271);
CN_in_sig(949)	<=	VN_out_sig(3272);
CN_in_sig(2117)	<=	VN_out_sig(3273);
CN_in_sig(2757)	<=	VN_out_sig(3274);
CN_in_sig(4421)	<=	VN_out_sig(3275);
CN_in_sig(957)	<=	VN_out_sig(3276);
CN_in_sig(2125)	<=	VN_out_sig(3277);
CN_in_sig(2765)	<=	VN_out_sig(3278);
CN_in_sig(4429)	<=	VN_out_sig(3279);
CN_in_sig(965)	<=	VN_out_sig(3280);
CN_in_sig(2133)	<=	VN_out_sig(3281);
CN_in_sig(2773)	<=	VN_out_sig(3282);
CN_in_sig(4437)	<=	VN_out_sig(3283);
CN_in_sig(973)	<=	VN_out_sig(3284);
CN_in_sig(2141)	<=	VN_out_sig(3285);
CN_in_sig(2781)	<=	VN_out_sig(3286);
CN_in_sig(4445)	<=	VN_out_sig(3287);
CN_in_sig(981)	<=	VN_out_sig(3288);
CN_in_sig(2149)	<=	VN_out_sig(3289);
CN_in_sig(2789)	<=	VN_out_sig(3290);
CN_in_sig(4453)	<=	VN_out_sig(3291);
CN_in_sig(989)	<=	VN_out_sig(3292);
CN_in_sig(2157)	<=	VN_out_sig(3293);
CN_in_sig(2797)	<=	VN_out_sig(3294);
CN_in_sig(4461)	<=	VN_out_sig(3295);
CN_in_sig(997)	<=	VN_out_sig(3296);
CN_in_sig(1733)	<=	VN_out_sig(3297);
CN_in_sig(2805)	<=	VN_out_sig(3298);
CN_in_sig(4469)	<=	VN_out_sig(3299);
CN_in_sig(1005)	<=	VN_out_sig(3300);
CN_in_sig(1741)	<=	VN_out_sig(3301);
CN_in_sig(2813)	<=	VN_out_sig(3302);
CN_in_sig(4477)	<=	VN_out_sig(3303);
CN_in_sig(1013)	<=	VN_out_sig(3304);
CN_in_sig(1749)	<=	VN_out_sig(3305);
CN_in_sig(2821)	<=	VN_out_sig(3306);
CN_in_sig(4485)	<=	VN_out_sig(3307);
CN_in_sig(1021)	<=	VN_out_sig(3308);
CN_in_sig(1757)	<=	VN_out_sig(3309);
CN_in_sig(2829)	<=	VN_out_sig(3310);
CN_in_sig(4493)	<=	VN_out_sig(3311);
CN_in_sig(1029)	<=	VN_out_sig(3312);
CN_in_sig(1765)	<=	VN_out_sig(3313);
CN_in_sig(2837)	<=	VN_out_sig(3314);
CN_in_sig(4501)	<=	VN_out_sig(3315);
CN_in_sig(1037)	<=	VN_out_sig(3316);
CN_in_sig(1773)	<=	VN_out_sig(3317);
CN_in_sig(2845)	<=	VN_out_sig(3318);
CN_in_sig(4509)	<=	VN_out_sig(3319);
CN_in_sig(1045)	<=	VN_out_sig(3320);
CN_in_sig(1781)	<=	VN_out_sig(3321);
CN_in_sig(2853)	<=	VN_out_sig(3322);
CN_in_sig(4517)	<=	VN_out_sig(3323);
CN_in_sig(1053)	<=	VN_out_sig(3324);
CN_in_sig(1789)	<=	VN_out_sig(3325);
CN_in_sig(2861)	<=	VN_out_sig(3326);
CN_in_sig(4525)	<=	VN_out_sig(3327);
CN_in_sig(1061)	<=	VN_out_sig(3328);
CN_in_sig(1797)	<=	VN_out_sig(3329);
CN_in_sig(2869)	<=	VN_out_sig(3330);
CN_in_sig(4533)	<=	VN_out_sig(3331);
CN_in_sig(1069)	<=	VN_out_sig(3332);
CN_in_sig(1805)	<=	VN_out_sig(3333);
CN_in_sig(2877)	<=	VN_out_sig(3334);
CN_in_sig(4541)	<=	VN_out_sig(3335);
CN_in_sig(1077)	<=	VN_out_sig(3336);
CN_in_sig(1813)	<=	VN_out_sig(3337);
CN_in_sig(2885)	<=	VN_out_sig(3338);
CN_in_sig(4549)	<=	VN_out_sig(3339);
CN_in_sig(1085)	<=	VN_out_sig(3340);
CN_in_sig(1821)	<=	VN_out_sig(3341);
CN_in_sig(2893)	<=	VN_out_sig(3342);
CN_in_sig(4557)	<=	VN_out_sig(3343);
CN_in_sig(1093)	<=	VN_out_sig(3344);
CN_in_sig(1829)	<=	VN_out_sig(3345);
CN_in_sig(2901)	<=	VN_out_sig(3346);
CN_in_sig(4565)	<=	VN_out_sig(3347);
CN_in_sig(1101)	<=	VN_out_sig(3348);
CN_in_sig(1837)	<=	VN_out_sig(3349);
CN_in_sig(2909)	<=	VN_out_sig(3350);
CN_in_sig(4573)	<=	VN_out_sig(3351);
CN_in_sig(1109)	<=	VN_out_sig(3352);
CN_in_sig(1845)	<=	VN_out_sig(3353);
CN_in_sig(2917)	<=	VN_out_sig(3354);
CN_in_sig(4581)	<=	VN_out_sig(3355);
CN_in_sig(1117)	<=	VN_out_sig(3356);
CN_in_sig(1853)	<=	VN_out_sig(3357);
CN_in_sig(2925)	<=	VN_out_sig(3358);
CN_in_sig(4589)	<=	VN_out_sig(3359);
CN_in_sig(1125)	<=	VN_out_sig(3360);
CN_in_sig(1861)	<=	VN_out_sig(3361);
CN_in_sig(2933)	<=	VN_out_sig(3362);
CN_in_sig(4597)	<=	VN_out_sig(3363);
CN_in_sig(1133)	<=	VN_out_sig(3364);
CN_in_sig(1869)	<=	VN_out_sig(3365);
CN_in_sig(2941)	<=	VN_out_sig(3366);
CN_in_sig(4605)	<=	VN_out_sig(3367);
CN_in_sig(1141)	<=	VN_out_sig(3368);
CN_in_sig(1877)	<=	VN_out_sig(3369);
CN_in_sig(2949)	<=	VN_out_sig(3370);
CN_in_sig(4613)	<=	VN_out_sig(3371);
CN_in_sig(1149)	<=	VN_out_sig(3372);
CN_in_sig(1885)	<=	VN_out_sig(3373);
CN_in_sig(2957)	<=	VN_out_sig(3374);
CN_in_sig(4621)	<=	VN_out_sig(3375);
CN_in_sig(1157)	<=	VN_out_sig(3376);
CN_in_sig(1893)	<=	VN_out_sig(3377);
CN_in_sig(2965)	<=	VN_out_sig(3378);
CN_in_sig(4629)	<=	VN_out_sig(3379);
CN_in_sig(1165)	<=	VN_out_sig(3380);
CN_in_sig(1901)	<=	VN_out_sig(3381);
CN_in_sig(2973)	<=	VN_out_sig(3382);
CN_in_sig(4637)	<=	VN_out_sig(3383);
CN_in_sig(1173)	<=	VN_out_sig(3384);
CN_in_sig(1909)	<=	VN_out_sig(3385);
CN_in_sig(2981)	<=	VN_out_sig(3386);
CN_in_sig(4645)	<=	VN_out_sig(3387);
CN_in_sig(1181)	<=	VN_out_sig(3388);
CN_in_sig(1917)	<=	VN_out_sig(3389);
CN_in_sig(2989)	<=	VN_out_sig(3390);
CN_in_sig(4653)	<=	VN_out_sig(3391);
CN_in_sig(1189)	<=	VN_out_sig(3392);
CN_in_sig(1925)	<=	VN_out_sig(3393);
CN_in_sig(2997)	<=	VN_out_sig(3394);
CN_in_sig(4661)	<=	VN_out_sig(3395);
CN_in_sig(1197)	<=	VN_out_sig(3396);
CN_in_sig(1933)	<=	VN_out_sig(3397);
CN_in_sig(3005)	<=	VN_out_sig(3398);
CN_in_sig(4669)	<=	VN_out_sig(3399);
CN_in_sig(1205)	<=	VN_out_sig(3400);
CN_in_sig(1941)	<=	VN_out_sig(3401);
CN_in_sig(3013)	<=	VN_out_sig(3402);
CN_in_sig(4677)	<=	VN_out_sig(3403);
CN_in_sig(1213)	<=	VN_out_sig(3404);
CN_in_sig(1949)	<=	VN_out_sig(3405);
CN_in_sig(3021)	<=	VN_out_sig(3406);
CN_in_sig(4685)	<=	VN_out_sig(3407);
CN_in_sig(1221)	<=	VN_out_sig(3408);
CN_in_sig(1957)	<=	VN_out_sig(3409);
CN_in_sig(2597)	<=	VN_out_sig(3410);
CN_in_sig(4693)	<=	VN_out_sig(3411);
CN_in_sig(1229)	<=	VN_out_sig(3412);
CN_in_sig(1965)	<=	VN_out_sig(3413);
CN_in_sig(2605)	<=	VN_out_sig(3414);
CN_in_sig(4701)	<=	VN_out_sig(3415);
CN_in_sig(1237)	<=	VN_out_sig(3416);
CN_in_sig(1973)	<=	VN_out_sig(3417);
CN_in_sig(2613)	<=	VN_out_sig(3418);
CN_in_sig(4709)	<=	VN_out_sig(3419);
CN_in_sig(1245)	<=	VN_out_sig(3420);
CN_in_sig(1981)	<=	VN_out_sig(3421);
CN_in_sig(2621)	<=	VN_out_sig(3422);
CN_in_sig(4717)	<=	VN_out_sig(3423);
CN_in_sig(1253)	<=	VN_out_sig(3424);
CN_in_sig(1989)	<=	VN_out_sig(3425);
CN_in_sig(2629)	<=	VN_out_sig(3426);
CN_in_sig(4725)	<=	VN_out_sig(3427);
CN_in_sig(1261)	<=	VN_out_sig(3428);
CN_in_sig(1997)	<=	VN_out_sig(3429);
CN_in_sig(2637)	<=	VN_out_sig(3430);
CN_in_sig(4733)	<=	VN_out_sig(3431);
CN_in_sig(1269)	<=	VN_out_sig(3432);
CN_in_sig(2005)	<=	VN_out_sig(3433);
CN_in_sig(2645)	<=	VN_out_sig(3434);
CN_in_sig(4741)	<=	VN_out_sig(3435);
CN_in_sig(1277)	<=	VN_out_sig(3436);
CN_in_sig(2013)	<=	VN_out_sig(3437);
CN_in_sig(2653)	<=	VN_out_sig(3438);
CN_in_sig(4749)	<=	VN_out_sig(3439);
CN_in_sig(1285)	<=	VN_out_sig(3440);
CN_in_sig(2021)	<=	VN_out_sig(3441);
CN_in_sig(2661)	<=	VN_out_sig(3442);
CN_in_sig(4325)	<=	VN_out_sig(3443);
CN_in_sig(1293)	<=	VN_out_sig(3444);
CN_in_sig(2029)	<=	VN_out_sig(3445);
CN_in_sig(2669)	<=	VN_out_sig(3446);
CN_in_sig(4333)	<=	VN_out_sig(3447);
CN_in_sig(869)	<=	VN_out_sig(3448);
CN_in_sig(2037)	<=	VN_out_sig(3449);
CN_in_sig(2677)	<=	VN_out_sig(3450);
CN_in_sig(4341)	<=	VN_out_sig(3451);
CN_in_sig(877)	<=	VN_out_sig(3452);
CN_in_sig(2045)	<=	VN_out_sig(3453);
CN_in_sig(2685)	<=	VN_out_sig(3454);
CN_in_sig(4349)	<=	VN_out_sig(3455);
CN_in_sig(85)	<=	VN_out_sig(3456);
CN_in_sig(1517)	<=	VN_out_sig(3457);
CN_in_sig(3853)	<=	VN_out_sig(3458);
CN_in_sig(5093)	<=	VN_out_sig(3459);
CN_in_sig(93)	<=	VN_out_sig(3460);
CN_in_sig(1525)	<=	VN_out_sig(3461);
CN_in_sig(3861)	<=	VN_out_sig(3462);
CN_in_sig(5101)	<=	VN_out_sig(3463);
CN_in_sig(101)	<=	VN_out_sig(3464);
CN_in_sig(1533)	<=	VN_out_sig(3465);
CN_in_sig(3869)	<=	VN_out_sig(3466);
CN_in_sig(5109)	<=	VN_out_sig(3467);
CN_in_sig(109)	<=	VN_out_sig(3468);
CN_in_sig(1541)	<=	VN_out_sig(3469);
CN_in_sig(3877)	<=	VN_out_sig(3470);
CN_in_sig(5117)	<=	VN_out_sig(3471);
CN_in_sig(117)	<=	VN_out_sig(3472);
CN_in_sig(1549)	<=	VN_out_sig(3473);
CN_in_sig(3885)	<=	VN_out_sig(3474);
CN_in_sig(5125)	<=	VN_out_sig(3475);
CN_in_sig(125)	<=	VN_out_sig(3476);
CN_in_sig(1557)	<=	VN_out_sig(3477);
CN_in_sig(3461)	<=	VN_out_sig(3478);
CN_in_sig(5133)	<=	VN_out_sig(3479);
CN_in_sig(133)	<=	VN_out_sig(3480);
CN_in_sig(1565)	<=	VN_out_sig(3481);
CN_in_sig(3469)	<=	VN_out_sig(3482);
CN_in_sig(5141)	<=	VN_out_sig(3483);
CN_in_sig(141)	<=	VN_out_sig(3484);
CN_in_sig(1573)	<=	VN_out_sig(3485);
CN_in_sig(3477)	<=	VN_out_sig(3486);
CN_in_sig(5149)	<=	VN_out_sig(3487);
CN_in_sig(149)	<=	VN_out_sig(3488);
CN_in_sig(1581)	<=	VN_out_sig(3489);
CN_in_sig(3485)	<=	VN_out_sig(3490);
CN_in_sig(5157)	<=	VN_out_sig(3491);
CN_in_sig(157)	<=	VN_out_sig(3492);
CN_in_sig(1589)	<=	VN_out_sig(3493);
CN_in_sig(3493)	<=	VN_out_sig(3494);
CN_in_sig(5165)	<=	VN_out_sig(3495);
CN_in_sig(165)	<=	VN_out_sig(3496);
CN_in_sig(1597)	<=	VN_out_sig(3497);
CN_in_sig(3501)	<=	VN_out_sig(3498);
CN_in_sig(5173)	<=	VN_out_sig(3499);
CN_in_sig(173)	<=	VN_out_sig(3500);
CN_in_sig(1605)	<=	VN_out_sig(3501);
CN_in_sig(3509)	<=	VN_out_sig(3502);
CN_in_sig(5181)	<=	VN_out_sig(3503);
CN_in_sig(181)	<=	VN_out_sig(3504);
CN_in_sig(1613)	<=	VN_out_sig(3505);
CN_in_sig(3517)	<=	VN_out_sig(3506);
CN_in_sig(4757)	<=	VN_out_sig(3507);
CN_in_sig(189)	<=	VN_out_sig(3508);
CN_in_sig(1621)	<=	VN_out_sig(3509);
CN_in_sig(3525)	<=	VN_out_sig(3510);
CN_in_sig(4765)	<=	VN_out_sig(3511);
CN_in_sig(197)	<=	VN_out_sig(3512);
CN_in_sig(1629)	<=	VN_out_sig(3513);
CN_in_sig(3533)	<=	VN_out_sig(3514);
CN_in_sig(4773)	<=	VN_out_sig(3515);
CN_in_sig(205)	<=	VN_out_sig(3516);
CN_in_sig(1637)	<=	VN_out_sig(3517);
CN_in_sig(3541)	<=	VN_out_sig(3518);
CN_in_sig(4781)	<=	VN_out_sig(3519);
CN_in_sig(213)	<=	VN_out_sig(3520);
CN_in_sig(1645)	<=	VN_out_sig(3521);
CN_in_sig(3549)	<=	VN_out_sig(3522);
CN_in_sig(4789)	<=	VN_out_sig(3523);
CN_in_sig(221)	<=	VN_out_sig(3524);
CN_in_sig(1653)	<=	VN_out_sig(3525);
CN_in_sig(3557)	<=	VN_out_sig(3526);
CN_in_sig(4797)	<=	VN_out_sig(3527);
CN_in_sig(229)	<=	VN_out_sig(3528);
CN_in_sig(1661)	<=	VN_out_sig(3529);
CN_in_sig(3565)	<=	VN_out_sig(3530);
CN_in_sig(4805)	<=	VN_out_sig(3531);
CN_in_sig(237)	<=	VN_out_sig(3532);
CN_in_sig(1669)	<=	VN_out_sig(3533);
CN_in_sig(3573)	<=	VN_out_sig(3534);
CN_in_sig(4813)	<=	VN_out_sig(3535);
CN_in_sig(245)	<=	VN_out_sig(3536);
CN_in_sig(1677)	<=	VN_out_sig(3537);
CN_in_sig(3581)	<=	VN_out_sig(3538);
CN_in_sig(4821)	<=	VN_out_sig(3539);
CN_in_sig(253)	<=	VN_out_sig(3540);
CN_in_sig(1685)	<=	VN_out_sig(3541);
CN_in_sig(3589)	<=	VN_out_sig(3542);
CN_in_sig(4829)	<=	VN_out_sig(3543);
CN_in_sig(261)	<=	VN_out_sig(3544);
CN_in_sig(1693)	<=	VN_out_sig(3545);
CN_in_sig(3597)	<=	VN_out_sig(3546);
CN_in_sig(4837)	<=	VN_out_sig(3547);
CN_in_sig(269)	<=	VN_out_sig(3548);
CN_in_sig(1701)	<=	VN_out_sig(3549);
CN_in_sig(3605)	<=	VN_out_sig(3550);
CN_in_sig(4845)	<=	VN_out_sig(3551);
CN_in_sig(277)	<=	VN_out_sig(3552);
CN_in_sig(1709)	<=	VN_out_sig(3553);
CN_in_sig(3613)	<=	VN_out_sig(3554);
CN_in_sig(4853)	<=	VN_out_sig(3555);
CN_in_sig(285)	<=	VN_out_sig(3556);
CN_in_sig(1717)	<=	VN_out_sig(3557);
CN_in_sig(3621)	<=	VN_out_sig(3558);
CN_in_sig(4861)	<=	VN_out_sig(3559);
CN_in_sig(293)	<=	VN_out_sig(3560);
CN_in_sig(1725)	<=	VN_out_sig(3561);
CN_in_sig(3629)	<=	VN_out_sig(3562);
CN_in_sig(4869)	<=	VN_out_sig(3563);
CN_in_sig(301)	<=	VN_out_sig(3564);
CN_in_sig(1301)	<=	VN_out_sig(3565);
CN_in_sig(3637)	<=	VN_out_sig(3566);
CN_in_sig(4877)	<=	VN_out_sig(3567);
CN_in_sig(309)	<=	VN_out_sig(3568);
CN_in_sig(1309)	<=	VN_out_sig(3569);
CN_in_sig(3645)	<=	VN_out_sig(3570);
CN_in_sig(4885)	<=	VN_out_sig(3571);
CN_in_sig(317)	<=	VN_out_sig(3572);
CN_in_sig(1317)	<=	VN_out_sig(3573);
CN_in_sig(3653)	<=	VN_out_sig(3574);
CN_in_sig(4893)	<=	VN_out_sig(3575);
CN_in_sig(325)	<=	VN_out_sig(3576);
CN_in_sig(1325)	<=	VN_out_sig(3577);
CN_in_sig(3661)	<=	VN_out_sig(3578);
CN_in_sig(4901)	<=	VN_out_sig(3579);
CN_in_sig(333)	<=	VN_out_sig(3580);
CN_in_sig(1333)	<=	VN_out_sig(3581);
CN_in_sig(3669)	<=	VN_out_sig(3582);
CN_in_sig(4909)	<=	VN_out_sig(3583);
CN_in_sig(341)	<=	VN_out_sig(3584);
CN_in_sig(1341)	<=	VN_out_sig(3585);
CN_in_sig(3677)	<=	VN_out_sig(3586);
CN_in_sig(4917)	<=	VN_out_sig(3587);
CN_in_sig(349)	<=	VN_out_sig(3588);
CN_in_sig(1349)	<=	VN_out_sig(3589);
CN_in_sig(3685)	<=	VN_out_sig(3590);
CN_in_sig(4925)	<=	VN_out_sig(3591);
CN_in_sig(357)	<=	VN_out_sig(3592);
CN_in_sig(1357)	<=	VN_out_sig(3593);
CN_in_sig(3693)	<=	VN_out_sig(3594);
CN_in_sig(4933)	<=	VN_out_sig(3595);
CN_in_sig(365)	<=	VN_out_sig(3596);
CN_in_sig(1365)	<=	VN_out_sig(3597);
CN_in_sig(3701)	<=	VN_out_sig(3598);
CN_in_sig(4941)	<=	VN_out_sig(3599);
CN_in_sig(373)	<=	VN_out_sig(3600);
CN_in_sig(1373)	<=	VN_out_sig(3601);
CN_in_sig(3709)	<=	VN_out_sig(3602);
CN_in_sig(4949)	<=	VN_out_sig(3603);
CN_in_sig(381)	<=	VN_out_sig(3604);
CN_in_sig(1381)	<=	VN_out_sig(3605);
CN_in_sig(3717)	<=	VN_out_sig(3606);
CN_in_sig(4957)	<=	VN_out_sig(3607);
CN_in_sig(389)	<=	VN_out_sig(3608);
CN_in_sig(1389)	<=	VN_out_sig(3609);
CN_in_sig(3725)	<=	VN_out_sig(3610);
CN_in_sig(4965)	<=	VN_out_sig(3611);
CN_in_sig(397)	<=	VN_out_sig(3612);
CN_in_sig(1397)	<=	VN_out_sig(3613);
CN_in_sig(3733)	<=	VN_out_sig(3614);
CN_in_sig(4973)	<=	VN_out_sig(3615);
CN_in_sig(405)	<=	VN_out_sig(3616);
CN_in_sig(1405)	<=	VN_out_sig(3617);
CN_in_sig(3741)	<=	VN_out_sig(3618);
CN_in_sig(4981)	<=	VN_out_sig(3619);
CN_in_sig(413)	<=	VN_out_sig(3620);
CN_in_sig(1413)	<=	VN_out_sig(3621);
CN_in_sig(3749)	<=	VN_out_sig(3622);
CN_in_sig(4989)	<=	VN_out_sig(3623);
CN_in_sig(421)	<=	VN_out_sig(3624);
CN_in_sig(1421)	<=	VN_out_sig(3625);
CN_in_sig(3757)	<=	VN_out_sig(3626);
CN_in_sig(4997)	<=	VN_out_sig(3627);
CN_in_sig(429)	<=	VN_out_sig(3628);
CN_in_sig(1429)	<=	VN_out_sig(3629);
CN_in_sig(3765)	<=	VN_out_sig(3630);
CN_in_sig(5005)	<=	VN_out_sig(3631);
CN_in_sig(5)	<=	VN_out_sig(3632);
CN_in_sig(1437)	<=	VN_out_sig(3633);
CN_in_sig(3773)	<=	VN_out_sig(3634);
CN_in_sig(5013)	<=	VN_out_sig(3635);
CN_in_sig(13)	<=	VN_out_sig(3636);
CN_in_sig(1445)	<=	VN_out_sig(3637);
CN_in_sig(3781)	<=	VN_out_sig(3638);
CN_in_sig(5021)	<=	VN_out_sig(3639);
CN_in_sig(21)	<=	VN_out_sig(3640);
CN_in_sig(1453)	<=	VN_out_sig(3641);
CN_in_sig(3789)	<=	VN_out_sig(3642);
CN_in_sig(5029)	<=	VN_out_sig(3643);
CN_in_sig(29)	<=	VN_out_sig(3644);
CN_in_sig(1461)	<=	VN_out_sig(3645);
CN_in_sig(3797)	<=	VN_out_sig(3646);
CN_in_sig(5037)	<=	VN_out_sig(3647);
CN_in_sig(37)	<=	VN_out_sig(3648);
CN_in_sig(1469)	<=	VN_out_sig(3649);
CN_in_sig(3805)	<=	VN_out_sig(3650);
CN_in_sig(5045)	<=	VN_out_sig(3651);
CN_in_sig(45)	<=	VN_out_sig(3652);
CN_in_sig(1477)	<=	VN_out_sig(3653);
CN_in_sig(3813)	<=	VN_out_sig(3654);
CN_in_sig(5053)	<=	VN_out_sig(3655);
CN_in_sig(53)	<=	VN_out_sig(3656);
CN_in_sig(1485)	<=	VN_out_sig(3657);
CN_in_sig(3821)	<=	VN_out_sig(3658);
CN_in_sig(5061)	<=	VN_out_sig(3659);
CN_in_sig(61)	<=	VN_out_sig(3660);
CN_in_sig(1493)	<=	VN_out_sig(3661);
CN_in_sig(3829)	<=	VN_out_sig(3662);
CN_in_sig(5069)	<=	VN_out_sig(3663);
CN_in_sig(69)	<=	VN_out_sig(3664);
CN_in_sig(1501)	<=	VN_out_sig(3665);
CN_in_sig(3837)	<=	VN_out_sig(3666);
CN_in_sig(5077)	<=	VN_out_sig(3667);
CN_in_sig(77)	<=	VN_out_sig(3668);
CN_in_sig(1509)	<=	VN_out_sig(3669);
CN_in_sig(3845)	<=	VN_out_sig(3670);
CN_in_sig(5085)	<=	VN_out_sig(3671);
CN_in_sig(597)	<=	VN_out_sig(3672);
CN_in_sig(2445)	<=	VN_out_sig(3673);
CN_in_sig(3237)	<=	VN_out_sig(3674);
CN_in_sig(4285)	<=	VN_out_sig(3675);
CN_in_sig(605)	<=	VN_out_sig(3676);
CN_in_sig(2453)	<=	VN_out_sig(3677);
CN_in_sig(3245)	<=	VN_out_sig(3678);
CN_in_sig(4293)	<=	VN_out_sig(3679);
CN_in_sig(613)	<=	VN_out_sig(3680);
CN_in_sig(2461)	<=	VN_out_sig(3681);
CN_in_sig(3253)	<=	VN_out_sig(3682);
CN_in_sig(4301)	<=	VN_out_sig(3683);
CN_in_sig(621)	<=	VN_out_sig(3684);
CN_in_sig(2469)	<=	VN_out_sig(3685);
CN_in_sig(3261)	<=	VN_out_sig(3686);
CN_in_sig(4309)	<=	VN_out_sig(3687);
CN_in_sig(629)	<=	VN_out_sig(3688);
CN_in_sig(2477)	<=	VN_out_sig(3689);
CN_in_sig(3269)	<=	VN_out_sig(3690);
CN_in_sig(4317)	<=	VN_out_sig(3691);
CN_in_sig(637)	<=	VN_out_sig(3692);
CN_in_sig(2485)	<=	VN_out_sig(3693);
CN_in_sig(3277)	<=	VN_out_sig(3694);
CN_in_sig(3893)	<=	VN_out_sig(3695);
CN_in_sig(645)	<=	VN_out_sig(3696);
CN_in_sig(2493)	<=	VN_out_sig(3697);
CN_in_sig(3285)	<=	VN_out_sig(3698);
CN_in_sig(3901)	<=	VN_out_sig(3699);
CN_in_sig(653)	<=	VN_out_sig(3700);
CN_in_sig(2501)	<=	VN_out_sig(3701);
CN_in_sig(3293)	<=	VN_out_sig(3702);
CN_in_sig(3909)	<=	VN_out_sig(3703);
CN_in_sig(661)	<=	VN_out_sig(3704);
CN_in_sig(2509)	<=	VN_out_sig(3705);
CN_in_sig(3301)	<=	VN_out_sig(3706);
CN_in_sig(3917)	<=	VN_out_sig(3707);
CN_in_sig(669)	<=	VN_out_sig(3708);
CN_in_sig(2517)	<=	VN_out_sig(3709);
CN_in_sig(3309)	<=	VN_out_sig(3710);
CN_in_sig(3925)	<=	VN_out_sig(3711);
CN_in_sig(677)	<=	VN_out_sig(3712);
CN_in_sig(2525)	<=	VN_out_sig(3713);
CN_in_sig(3317)	<=	VN_out_sig(3714);
CN_in_sig(3933)	<=	VN_out_sig(3715);
CN_in_sig(685)	<=	VN_out_sig(3716);
CN_in_sig(2533)	<=	VN_out_sig(3717);
CN_in_sig(3325)	<=	VN_out_sig(3718);
CN_in_sig(3941)	<=	VN_out_sig(3719);
CN_in_sig(693)	<=	VN_out_sig(3720);
CN_in_sig(2541)	<=	VN_out_sig(3721);
CN_in_sig(3333)	<=	VN_out_sig(3722);
CN_in_sig(3949)	<=	VN_out_sig(3723);
CN_in_sig(701)	<=	VN_out_sig(3724);
CN_in_sig(2549)	<=	VN_out_sig(3725);
CN_in_sig(3341)	<=	VN_out_sig(3726);
CN_in_sig(3957)	<=	VN_out_sig(3727);
CN_in_sig(709)	<=	VN_out_sig(3728);
CN_in_sig(2557)	<=	VN_out_sig(3729);
CN_in_sig(3349)	<=	VN_out_sig(3730);
CN_in_sig(3965)	<=	VN_out_sig(3731);
CN_in_sig(717)	<=	VN_out_sig(3732);
CN_in_sig(2565)	<=	VN_out_sig(3733);
CN_in_sig(3357)	<=	VN_out_sig(3734);
CN_in_sig(3973)	<=	VN_out_sig(3735);
CN_in_sig(725)	<=	VN_out_sig(3736);
CN_in_sig(2573)	<=	VN_out_sig(3737);
CN_in_sig(3365)	<=	VN_out_sig(3738);
CN_in_sig(3981)	<=	VN_out_sig(3739);
CN_in_sig(733)	<=	VN_out_sig(3740);
CN_in_sig(2581)	<=	VN_out_sig(3741);
CN_in_sig(3373)	<=	VN_out_sig(3742);
CN_in_sig(3989)	<=	VN_out_sig(3743);
CN_in_sig(741)	<=	VN_out_sig(3744);
CN_in_sig(2589)	<=	VN_out_sig(3745);
CN_in_sig(3381)	<=	VN_out_sig(3746);
CN_in_sig(3997)	<=	VN_out_sig(3747);
CN_in_sig(749)	<=	VN_out_sig(3748);
CN_in_sig(2165)	<=	VN_out_sig(3749);
CN_in_sig(3389)	<=	VN_out_sig(3750);
CN_in_sig(4005)	<=	VN_out_sig(3751);
CN_in_sig(757)	<=	VN_out_sig(3752);
CN_in_sig(2173)	<=	VN_out_sig(3753);
CN_in_sig(3397)	<=	VN_out_sig(3754);
CN_in_sig(4013)	<=	VN_out_sig(3755);
CN_in_sig(765)	<=	VN_out_sig(3756);
CN_in_sig(2181)	<=	VN_out_sig(3757);
CN_in_sig(3405)	<=	VN_out_sig(3758);
CN_in_sig(4021)	<=	VN_out_sig(3759);
CN_in_sig(773)	<=	VN_out_sig(3760);
CN_in_sig(2189)	<=	VN_out_sig(3761);
CN_in_sig(3413)	<=	VN_out_sig(3762);
CN_in_sig(4029)	<=	VN_out_sig(3763);
CN_in_sig(781)	<=	VN_out_sig(3764);
CN_in_sig(2197)	<=	VN_out_sig(3765);
CN_in_sig(3421)	<=	VN_out_sig(3766);
CN_in_sig(4037)	<=	VN_out_sig(3767);
CN_in_sig(789)	<=	VN_out_sig(3768);
CN_in_sig(2205)	<=	VN_out_sig(3769);
CN_in_sig(3429)	<=	VN_out_sig(3770);
CN_in_sig(4045)	<=	VN_out_sig(3771);
CN_in_sig(797)	<=	VN_out_sig(3772);
CN_in_sig(2213)	<=	VN_out_sig(3773);
CN_in_sig(3437)	<=	VN_out_sig(3774);
CN_in_sig(4053)	<=	VN_out_sig(3775);
CN_in_sig(805)	<=	VN_out_sig(3776);
CN_in_sig(2221)	<=	VN_out_sig(3777);
CN_in_sig(3445)	<=	VN_out_sig(3778);
CN_in_sig(4061)	<=	VN_out_sig(3779);
CN_in_sig(813)	<=	VN_out_sig(3780);
CN_in_sig(2229)	<=	VN_out_sig(3781);
CN_in_sig(3453)	<=	VN_out_sig(3782);
CN_in_sig(4069)	<=	VN_out_sig(3783);
CN_in_sig(821)	<=	VN_out_sig(3784);
CN_in_sig(2237)	<=	VN_out_sig(3785);
CN_in_sig(3029)	<=	VN_out_sig(3786);
CN_in_sig(4077)	<=	VN_out_sig(3787);
CN_in_sig(829)	<=	VN_out_sig(3788);
CN_in_sig(2245)	<=	VN_out_sig(3789);
CN_in_sig(3037)	<=	VN_out_sig(3790);
CN_in_sig(4085)	<=	VN_out_sig(3791);
CN_in_sig(837)	<=	VN_out_sig(3792);
CN_in_sig(2253)	<=	VN_out_sig(3793);
CN_in_sig(3045)	<=	VN_out_sig(3794);
CN_in_sig(4093)	<=	VN_out_sig(3795);
CN_in_sig(845)	<=	VN_out_sig(3796);
CN_in_sig(2261)	<=	VN_out_sig(3797);
CN_in_sig(3053)	<=	VN_out_sig(3798);
CN_in_sig(4101)	<=	VN_out_sig(3799);
CN_in_sig(853)	<=	VN_out_sig(3800);
CN_in_sig(2269)	<=	VN_out_sig(3801);
CN_in_sig(3061)	<=	VN_out_sig(3802);
CN_in_sig(4109)	<=	VN_out_sig(3803);
CN_in_sig(861)	<=	VN_out_sig(3804);
CN_in_sig(2277)	<=	VN_out_sig(3805);
CN_in_sig(3069)	<=	VN_out_sig(3806);
CN_in_sig(4117)	<=	VN_out_sig(3807);
CN_in_sig(437)	<=	VN_out_sig(3808);
CN_in_sig(2285)	<=	VN_out_sig(3809);
CN_in_sig(3077)	<=	VN_out_sig(3810);
CN_in_sig(4125)	<=	VN_out_sig(3811);
CN_in_sig(445)	<=	VN_out_sig(3812);
CN_in_sig(2293)	<=	VN_out_sig(3813);
CN_in_sig(3085)	<=	VN_out_sig(3814);
CN_in_sig(4133)	<=	VN_out_sig(3815);
CN_in_sig(453)	<=	VN_out_sig(3816);
CN_in_sig(2301)	<=	VN_out_sig(3817);
CN_in_sig(3093)	<=	VN_out_sig(3818);
CN_in_sig(4141)	<=	VN_out_sig(3819);
CN_in_sig(461)	<=	VN_out_sig(3820);
CN_in_sig(2309)	<=	VN_out_sig(3821);
CN_in_sig(3101)	<=	VN_out_sig(3822);
CN_in_sig(4149)	<=	VN_out_sig(3823);
CN_in_sig(469)	<=	VN_out_sig(3824);
CN_in_sig(2317)	<=	VN_out_sig(3825);
CN_in_sig(3109)	<=	VN_out_sig(3826);
CN_in_sig(4157)	<=	VN_out_sig(3827);
CN_in_sig(477)	<=	VN_out_sig(3828);
CN_in_sig(2325)	<=	VN_out_sig(3829);
CN_in_sig(3117)	<=	VN_out_sig(3830);
CN_in_sig(4165)	<=	VN_out_sig(3831);
CN_in_sig(485)	<=	VN_out_sig(3832);
CN_in_sig(2333)	<=	VN_out_sig(3833);
CN_in_sig(3125)	<=	VN_out_sig(3834);
CN_in_sig(4173)	<=	VN_out_sig(3835);
CN_in_sig(493)	<=	VN_out_sig(3836);
CN_in_sig(2341)	<=	VN_out_sig(3837);
CN_in_sig(3133)	<=	VN_out_sig(3838);
CN_in_sig(4181)	<=	VN_out_sig(3839);
CN_in_sig(501)	<=	VN_out_sig(3840);
CN_in_sig(2349)	<=	VN_out_sig(3841);
CN_in_sig(3141)	<=	VN_out_sig(3842);
CN_in_sig(4189)	<=	VN_out_sig(3843);
CN_in_sig(509)	<=	VN_out_sig(3844);
CN_in_sig(2357)	<=	VN_out_sig(3845);
CN_in_sig(3149)	<=	VN_out_sig(3846);
CN_in_sig(4197)	<=	VN_out_sig(3847);
CN_in_sig(517)	<=	VN_out_sig(3848);
CN_in_sig(2365)	<=	VN_out_sig(3849);
CN_in_sig(3157)	<=	VN_out_sig(3850);
CN_in_sig(4205)	<=	VN_out_sig(3851);
CN_in_sig(525)	<=	VN_out_sig(3852);
CN_in_sig(2373)	<=	VN_out_sig(3853);
CN_in_sig(3165)	<=	VN_out_sig(3854);
CN_in_sig(4213)	<=	VN_out_sig(3855);
CN_in_sig(533)	<=	VN_out_sig(3856);
CN_in_sig(2381)	<=	VN_out_sig(3857);
CN_in_sig(3173)	<=	VN_out_sig(3858);
CN_in_sig(4221)	<=	VN_out_sig(3859);
CN_in_sig(541)	<=	VN_out_sig(3860);
CN_in_sig(2389)	<=	VN_out_sig(3861);
CN_in_sig(3181)	<=	VN_out_sig(3862);
CN_in_sig(4229)	<=	VN_out_sig(3863);
CN_in_sig(549)	<=	VN_out_sig(3864);
CN_in_sig(2397)	<=	VN_out_sig(3865);
CN_in_sig(3189)	<=	VN_out_sig(3866);
CN_in_sig(4237)	<=	VN_out_sig(3867);
CN_in_sig(557)	<=	VN_out_sig(3868);
CN_in_sig(2405)	<=	VN_out_sig(3869);
CN_in_sig(3197)	<=	VN_out_sig(3870);
CN_in_sig(4245)	<=	VN_out_sig(3871);
CN_in_sig(565)	<=	VN_out_sig(3872);
CN_in_sig(2413)	<=	VN_out_sig(3873);
CN_in_sig(3205)	<=	VN_out_sig(3874);
CN_in_sig(4253)	<=	VN_out_sig(3875);
CN_in_sig(573)	<=	VN_out_sig(3876);
CN_in_sig(2421)	<=	VN_out_sig(3877);
CN_in_sig(3213)	<=	VN_out_sig(3878);
CN_in_sig(4261)	<=	VN_out_sig(3879);
CN_in_sig(581)	<=	VN_out_sig(3880);
CN_in_sig(2429)	<=	VN_out_sig(3881);
CN_in_sig(3221)	<=	VN_out_sig(3882);
CN_in_sig(4269)	<=	VN_out_sig(3883);
CN_in_sig(589)	<=	VN_out_sig(3884);
CN_in_sig(2437)	<=	VN_out_sig(3885);
CN_in_sig(3229)	<=	VN_out_sig(3886);
CN_in_sig(4277)	<=	VN_out_sig(3887);
CN_in_sig(374)	<=	VN_out_sig(3888);
CN_in_sig(1702)	<=	VN_out_sig(3889);
CN_in_sig(3694)	<=	VN_out_sig(3890);
CN_in_sig(5126)	<=	VN_out_sig(3891);
CN_in_sig(382)	<=	VN_out_sig(3892);
CN_in_sig(1710)	<=	VN_out_sig(3893);
CN_in_sig(3702)	<=	VN_out_sig(3894);
CN_in_sig(5134)	<=	VN_out_sig(3895);
CN_in_sig(390)	<=	VN_out_sig(3896);
CN_in_sig(1718)	<=	VN_out_sig(3897);
CN_in_sig(3710)	<=	VN_out_sig(3898);
CN_in_sig(5142)	<=	VN_out_sig(3899);
CN_in_sig(398)	<=	VN_out_sig(3900);
CN_in_sig(1726)	<=	VN_out_sig(3901);
CN_in_sig(3718)	<=	VN_out_sig(3902);
CN_in_sig(5150)	<=	VN_out_sig(3903);
CN_in_sig(406)	<=	VN_out_sig(3904);
CN_in_sig(1302)	<=	VN_out_sig(3905);
CN_in_sig(3726)	<=	VN_out_sig(3906);
CN_in_sig(5158)	<=	VN_out_sig(3907);
CN_in_sig(414)	<=	VN_out_sig(3908);
CN_in_sig(1310)	<=	VN_out_sig(3909);
CN_in_sig(3734)	<=	VN_out_sig(3910);
CN_in_sig(5166)	<=	VN_out_sig(3911);
CN_in_sig(422)	<=	VN_out_sig(3912);
CN_in_sig(1318)	<=	VN_out_sig(3913);
CN_in_sig(3742)	<=	VN_out_sig(3914);
CN_in_sig(5174)	<=	VN_out_sig(3915);
CN_in_sig(430)	<=	VN_out_sig(3916);
CN_in_sig(1326)	<=	VN_out_sig(3917);
CN_in_sig(3750)	<=	VN_out_sig(3918);
CN_in_sig(5182)	<=	VN_out_sig(3919);
CN_in_sig(6)	<=	VN_out_sig(3920);
CN_in_sig(1334)	<=	VN_out_sig(3921);
CN_in_sig(3758)	<=	VN_out_sig(3922);
CN_in_sig(4758)	<=	VN_out_sig(3923);
CN_in_sig(14)	<=	VN_out_sig(3924);
CN_in_sig(1342)	<=	VN_out_sig(3925);
CN_in_sig(3766)	<=	VN_out_sig(3926);
CN_in_sig(4766)	<=	VN_out_sig(3927);
CN_in_sig(22)	<=	VN_out_sig(3928);
CN_in_sig(1350)	<=	VN_out_sig(3929);
CN_in_sig(3774)	<=	VN_out_sig(3930);
CN_in_sig(4774)	<=	VN_out_sig(3931);
CN_in_sig(30)	<=	VN_out_sig(3932);
CN_in_sig(1358)	<=	VN_out_sig(3933);
CN_in_sig(3782)	<=	VN_out_sig(3934);
CN_in_sig(4782)	<=	VN_out_sig(3935);
CN_in_sig(38)	<=	VN_out_sig(3936);
CN_in_sig(1366)	<=	VN_out_sig(3937);
CN_in_sig(3790)	<=	VN_out_sig(3938);
CN_in_sig(4790)	<=	VN_out_sig(3939);
CN_in_sig(46)	<=	VN_out_sig(3940);
CN_in_sig(1374)	<=	VN_out_sig(3941);
CN_in_sig(3798)	<=	VN_out_sig(3942);
CN_in_sig(4798)	<=	VN_out_sig(3943);
CN_in_sig(54)	<=	VN_out_sig(3944);
CN_in_sig(1382)	<=	VN_out_sig(3945);
CN_in_sig(3806)	<=	VN_out_sig(3946);
CN_in_sig(4806)	<=	VN_out_sig(3947);
CN_in_sig(62)	<=	VN_out_sig(3948);
CN_in_sig(1390)	<=	VN_out_sig(3949);
CN_in_sig(3814)	<=	VN_out_sig(3950);
CN_in_sig(4814)	<=	VN_out_sig(3951);
CN_in_sig(70)	<=	VN_out_sig(3952);
CN_in_sig(1398)	<=	VN_out_sig(3953);
CN_in_sig(3822)	<=	VN_out_sig(3954);
CN_in_sig(4822)	<=	VN_out_sig(3955);
CN_in_sig(78)	<=	VN_out_sig(3956);
CN_in_sig(1406)	<=	VN_out_sig(3957);
CN_in_sig(3830)	<=	VN_out_sig(3958);
CN_in_sig(4830)	<=	VN_out_sig(3959);
CN_in_sig(86)	<=	VN_out_sig(3960);
CN_in_sig(1414)	<=	VN_out_sig(3961);
CN_in_sig(3838)	<=	VN_out_sig(3962);
CN_in_sig(4838)	<=	VN_out_sig(3963);
CN_in_sig(94)	<=	VN_out_sig(3964);
CN_in_sig(1422)	<=	VN_out_sig(3965);
CN_in_sig(3846)	<=	VN_out_sig(3966);
CN_in_sig(4846)	<=	VN_out_sig(3967);
CN_in_sig(102)	<=	VN_out_sig(3968);
CN_in_sig(1430)	<=	VN_out_sig(3969);
CN_in_sig(3854)	<=	VN_out_sig(3970);
CN_in_sig(4854)	<=	VN_out_sig(3971);
CN_in_sig(110)	<=	VN_out_sig(3972);
CN_in_sig(1438)	<=	VN_out_sig(3973);
CN_in_sig(3862)	<=	VN_out_sig(3974);
CN_in_sig(4862)	<=	VN_out_sig(3975);
CN_in_sig(118)	<=	VN_out_sig(3976);
CN_in_sig(1446)	<=	VN_out_sig(3977);
CN_in_sig(3870)	<=	VN_out_sig(3978);
CN_in_sig(4870)	<=	VN_out_sig(3979);
CN_in_sig(126)	<=	VN_out_sig(3980);
CN_in_sig(1454)	<=	VN_out_sig(3981);
CN_in_sig(3878)	<=	VN_out_sig(3982);
CN_in_sig(4878)	<=	VN_out_sig(3983);
CN_in_sig(134)	<=	VN_out_sig(3984);
CN_in_sig(1462)	<=	VN_out_sig(3985);
CN_in_sig(3886)	<=	VN_out_sig(3986);
CN_in_sig(4886)	<=	VN_out_sig(3987);
CN_in_sig(142)	<=	VN_out_sig(3988);
CN_in_sig(1470)	<=	VN_out_sig(3989);
CN_in_sig(3462)	<=	VN_out_sig(3990);
CN_in_sig(4894)	<=	VN_out_sig(3991);
CN_in_sig(150)	<=	VN_out_sig(3992);
CN_in_sig(1478)	<=	VN_out_sig(3993);
CN_in_sig(3470)	<=	VN_out_sig(3994);
CN_in_sig(4902)	<=	VN_out_sig(3995);
CN_in_sig(158)	<=	VN_out_sig(3996);
CN_in_sig(1486)	<=	VN_out_sig(3997);
CN_in_sig(3478)	<=	VN_out_sig(3998);
CN_in_sig(4910)	<=	VN_out_sig(3999);
CN_in_sig(166)	<=	VN_out_sig(4000);
CN_in_sig(1494)	<=	VN_out_sig(4001);
CN_in_sig(3486)	<=	VN_out_sig(4002);
CN_in_sig(4918)	<=	VN_out_sig(4003);
CN_in_sig(174)	<=	VN_out_sig(4004);
CN_in_sig(1502)	<=	VN_out_sig(4005);
CN_in_sig(3494)	<=	VN_out_sig(4006);
CN_in_sig(4926)	<=	VN_out_sig(4007);
CN_in_sig(182)	<=	VN_out_sig(4008);
CN_in_sig(1510)	<=	VN_out_sig(4009);
CN_in_sig(3502)	<=	VN_out_sig(4010);
CN_in_sig(4934)	<=	VN_out_sig(4011);
CN_in_sig(190)	<=	VN_out_sig(4012);
CN_in_sig(1518)	<=	VN_out_sig(4013);
CN_in_sig(3510)	<=	VN_out_sig(4014);
CN_in_sig(4942)	<=	VN_out_sig(4015);
CN_in_sig(198)	<=	VN_out_sig(4016);
CN_in_sig(1526)	<=	VN_out_sig(4017);
CN_in_sig(3518)	<=	VN_out_sig(4018);
CN_in_sig(4950)	<=	VN_out_sig(4019);
CN_in_sig(206)	<=	VN_out_sig(4020);
CN_in_sig(1534)	<=	VN_out_sig(4021);
CN_in_sig(3526)	<=	VN_out_sig(4022);
CN_in_sig(4958)	<=	VN_out_sig(4023);
CN_in_sig(214)	<=	VN_out_sig(4024);
CN_in_sig(1542)	<=	VN_out_sig(4025);
CN_in_sig(3534)	<=	VN_out_sig(4026);
CN_in_sig(4966)	<=	VN_out_sig(4027);
CN_in_sig(222)	<=	VN_out_sig(4028);
CN_in_sig(1550)	<=	VN_out_sig(4029);
CN_in_sig(3542)	<=	VN_out_sig(4030);
CN_in_sig(4974)	<=	VN_out_sig(4031);
CN_in_sig(230)	<=	VN_out_sig(4032);
CN_in_sig(1558)	<=	VN_out_sig(4033);
CN_in_sig(3550)	<=	VN_out_sig(4034);
CN_in_sig(4982)	<=	VN_out_sig(4035);
CN_in_sig(238)	<=	VN_out_sig(4036);
CN_in_sig(1566)	<=	VN_out_sig(4037);
CN_in_sig(3558)	<=	VN_out_sig(4038);
CN_in_sig(4990)	<=	VN_out_sig(4039);
CN_in_sig(246)	<=	VN_out_sig(4040);
CN_in_sig(1574)	<=	VN_out_sig(4041);
CN_in_sig(3566)	<=	VN_out_sig(4042);
CN_in_sig(4998)	<=	VN_out_sig(4043);
CN_in_sig(254)	<=	VN_out_sig(4044);
CN_in_sig(1582)	<=	VN_out_sig(4045);
CN_in_sig(3574)	<=	VN_out_sig(4046);
CN_in_sig(5006)	<=	VN_out_sig(4047);
CN_in_sig(262)	<=	VN_out_sig(4048);
CN_in_sig(1590)	<=	VN_out_sig(4049);
CN_in_sig(3582)	<=	VN_out_sig(4050);
CN_in_sig(5014)	<=	VN_out_sig(4051);
CN_in_sig(270)	<=	VN_out_sig(4052);
CN_in_sig(1598)	<=	VN_out_sig(4053);
CN_in_sig(3590)	<=	VN_out_sig(4054);
CN_in_sig(5022)	<=	VN_out_sig(4055);
CN_in_sig(278)	<=	VN_out_sig(4056);
CN_in_sig(1606)	<=	VN_out_sig(4057);
CN_in_sig(3598)	<=	VN_out_sig(4058);
CN_in_sig(5030)	<=	VN_out_sig(4059);
CN_in_sig(286)	<=	VN_out_sig(4060);
CN_in_sig(1614)	<=	VN_out_sig(4061);
CN_in_sig(3606)	<=	VN_out_sig(4062);
CN_in_sig(5038)	<=	VN_out_sig(4063);
CN_in_sig(294)	<=	VN_out_sig(4064);
CN_in_sig(1622)	<=	VN_out_sig(4065);
CN_in_sig(3614)	<=	VN_out_sig(4066);
CN_in_sig(5046)	<=	VN_out_sig(4067);
CN_in_sig(302)	<=	VN_out_sig(4068);
CN_in_sig(1630)	<=	VN_out_sig(4069);
CN_in_sig(3622)	<=	VN_out_sig(4070);
CN_in_sig(5054)	<=	VN_out_sig(4071);
CN_in_sig(310)	<=	VN_out_sig(4072);
CN_in_sig(1638)	<=	VN_out_sig(4073);
CN_in_sig(3630)	<=	VN_out_sig(4074);
CN_in_sig(5062)	<=	VN_out_sig(4075);
CN_in_sig(318)	<=	VN_out_sig(4076);
CN_in_sig(1646)	<=	VN_out_sig(4077);
CN_in_sig(3638)	<=	VN_out_sig(4078);
CN_in_sig(5070)	<=	VN_out_sig(4079);
CN_in_sig(326)	<=	VN_out_sig(4080);
CN_in_sig(1654)	<=	VN_out_sig(4081);
CN_in_sig(3646)	<=	VN_out_sig(4082);
CN_in_sig(5078)	<=	VN_out_sig(4083);
CN_in_sig(334)	<=	VN_out_sig(4084);
CN_in_sig(1662)	<=	VN_out_sig(4085);
CN_in_sig(3654)	<=	VN_out_sig(4086);
CN_in_sig(5086)	<=	VN_out_sig(4087);
CN_in_sig(342)	<=	VN_out_sig(4088);
CN_in_sig(1670)	<=	VN_out_sig(4089);
CN_in_sig(3662)	<=	VN_out_sig(4090);
CN_in_sig(5094)	<=	VN_out_sig(4091);
CN_in_sig(350)	<=	VN_out_sig(4092);
CN_in_sig(1678)	<=	VN_out_sig(4093);
CN_in_sig(3670)	<=	VN_out_sig(4094);
CN_in_sig(5102)	<=	VN_out_sig(4095);
CN_in_sig(358)	<=	VN_out_sig(4096);
CN_in_sig(1686)	<=	VN_out_sig(4097);
CN_in_sig(3678)	<=	VN_out_sig(4098);
CN_in_sig(5110)	<=	VN_out_sig(4099);
CN_in_sig(366)	<=	VN_out_sig(4100);
CN_in_sig(1694)	<=	VN_out_sig(4101);
CN_in_sig(3686)	<=	VN_out_sig(4102);
CN_in_sig(5118)	<=	VN_out_sig(4103);
CN_in_sig(750)	<=	VN_out_sig(4104);
CN_in_sig(2294)	<=	VN_out_sig(4105);
CN_in_sig(2694)	<=	VN_out_sig(4106);
CN_in_sig(4046)	<=	VN_out_sig(4107);
CN_in_sig(758)	<=	VN_out_sig(4108);
CN_in_sig(2302)	<=	VN_out_sig(4109);
CN_in_sig(2702)	<=	VN_out_sig(4110);
CN_in_sig(4054)	<=	VN_out_sig(4111);
CN_in_sig(766)	<=	VN_out_sig(4112);
CN_in_sig(2310)	<=	VN_out_sig(4113);
CN_in_sig(2710)	<=	VN_out_sig(4114);
CN_in_sig(4062)	<=	VN_out_sig(4115);
CN_in_sig(774)	<=	VN_out_sig(4116);
CN_in_sig(2318)	<=	VN_out_sig(4117);
CN_in_sig(2718)	<=	VN_out_sig(4118);
CN_in_sig(4070)	<=	VN_out_sig(4119);
CN_in_sig(782)	<=	VN_out_sig(4120);
CN_in_sig(2326)	<=	VN_out_sig(4121);
CN_in_sig(2726)	<=	VN_out_sig(4122);
CN_in_sig(4078)	<=	VN_out_sig(4123);
CN_in_sig(790)	<=	VN_out_sig(4124);
CN_in_sig(2334)	<=	VN_out_sig(4125);
CN_in_sig(2734)	<=	VN_out_sig(4126);
CN_in_sig(4086)	<=	VN_out_sig(4127);
CN_in_sig(798)	<=	VN_out_sig(4128);
CN_in_sig(2342)	<=	VN_out_sig(4129);
CN_in_sig(2742)	<=	VN_out_sig(4130);
CN_in_sig(4094)	<=	VN_out_sig(4131);
CN_in_sig(806)	<=	VN_out_sig(4132);
CN_in_sig(2350)	<=	VN_out_sig(4133);
CN_in_sig(2750)	<=	VN_out_sig(4134);
CN_in_sig(4102)	<=	VN_out_sig(4135);
CN_in_sig(814)	<=	VN_out_sig(4136);
CN_in_sig(2358)	<=	VN_out_sig(4137);
CN_in_sig(2758)	<=	VN_out_sig(4138);
CN_in_sig(4110)	<=	VN_out_sig(4139);
CN_in_sig(822)	<=	VN_out_sig(4140);
CN_in_sig(2366)	<=	VN_out_sig(4141);
CN_in_sig(2766)	<=	VN_out_sig(4142);
CN_in_sig(4118)	<=	VN_out_sig(4143);
CN_in_sig(830)	<=	VN_out_sig(4144);
CN_in_sig(2374)	<=	VN_out_sig(4145);
CN_in_sig(2774)	<=	VN_out_sig(4146);
CN_in_sig(4126)	<=	VN_out_sig(4147);
CN_in_sig(838)	<=	VN_out_sig(4148);
CN_in_sig(2382)	<=	VN_out_sig(4149);
CN_in_sig(2782)	<=	VN_out_sig(4150);
CN_in_sig(4134)	<=	VN_out_sig(4151);
CN_in_sig(846)	<=	VN_out_sig(4152);
CN_in_sig(2390)	<=	VN_out_sig(4153);
CN_in_sig(2790)	<=	VN_out_sig(4154);
CN_in_sig(4142)	<=	VN_out_sig(4155);
CN_in_sig(854)	<=	VN_out_sig(4156);
CN_in_sig(2398)	<=	VN_out_sig(4157);
CN_in_sig(2798)	<=	VN_out_sig(4158);
CN_in_sig(4150)	<=	VN_out_sig(4159);
CN_in_sig(862)	<=	VN_out_sig(4160);
CN_in_sig(2406)	<=	VN_out_sig(4161);
CN_in_sig(2806)	<=	VN_out_sig(4162);
CN_in_sig(4158)	<=	VN_out_sig(4163);
CN_in_sig(438)	<=	VN_out_sig(4164);
CN_in_sig(2414)	<=	VN_out_sig(4165);
CN_in_sig(2814)	<=	VN_out_sig(4166);
CN_in_sig(4166)	<=	VN_out_sig(4167);
CN_in_sig(446)	<=	VN_out_sig(4168);
CN_in_sig(2422)	<=	VN_out_sig(4169);
CN_in_sig(2822)	<=	VN_out_sig(4170);
CN_in_sig(4174)	<=	VN_out_sig(4171);
CN_in_sig(454)	<=	VN_out_sig(4172);
CN_in_sig(2430)	<=	VN_out_sig(4173);
CN_in_sig(2830)	<=	VN_out_sig(4174);
CN_in_sig(4182)	<=	VN_out_sig(4175);
CN_in_sig(462)	<=	VN_out_sig(4176);
CN_in_sig(2438)	<=	VN_out_sig(4177);
CN_in_sig(2838)	<=	VN_out_sig(4178);
CN_in_sig(4190)	<=	VN_out_sig(4179);
CN_in_sig(470)	<=	VN_out_sig(4180);
CN_in_sig(2446)	<=	VN_out_sig(4181);
CN_in_sig(2846)	<=	VN_out_sig(4182);
CN_in_sig(4198)	<=	VN_out_sig(4183);
CN_in_sig(478)	<=	VN_out_sig(4184);
CN_in_sig(2454)	<=	VN_out_sig(4185);
CN_in_sig(2854)	<=	VN_out_sig(4186);
CN_in_sig(4206)	<=	VN_out_sig(4187);
CN_in_sig(486)	<=	VN_out_sig(4188);
CN_in_sig(2462)	<=	VN_out_sig(4189);
CN_in_sig(2862)	<=	VN_out_sig(4190);
CN_in_sig(4214)	<=	VN_out_sig(4191);
CN_in_sig(494)	<=	VN_out_sig(4192);
CN_in_sig(2470)	<=	VN_out_sig(4193);
CN_in_sig(2870)	<=	VN_out_sig(4194);
CN_in_sig(4222)	<=	VN_out_sig(4195);
CN_in_sig(502)	<=	VN_out_sig(4196);
CN_in_sig(2478)	<=	VN_out_sig(4197);
CN_in_sig(2878)	<=	VN_out_sig(4198);
CN_in_sig(4230)	<=	VN_out_sig(4199);
CN_in_sig(510)	<=	VN_out_sig(4200);
CN_in_sig(2486)	<=	VN_out_sig(4201);
CN_in_sig(2886)	<=	VN_out_sig(4202);
CN_in_sig(4238)	<=	VN_out_sig(4203);
CN_in_sig(518)	<=	VN_out_sig(4204);
CN_in_sig(2494)	<=	VN_out_sig(4205);
CN_in_sig(2894)	<=	VN_out_sig(4206);
CN_in_sig(4246)	<=	VN_out_sig(4207);
CN_in_sig(526)	<=	VN_out_sig(4208);
CN_in_sig(2502)	<=	VN_out_sig(4209);
CN_in_sig(2902)	<=	VN_out_sig(4210);
CN_in_sig(4254)	<=	VN_out_sig(4211);
CN_in_sig(534)	<=	VN_out_sig(4212);
CN_in_sig(2510)	<=	VN_out_sig(4213);
CN_in_sig(2910)	<=	VN_out_sig(4214);
CN_in_sig(4262)	<=	VN_out_sig(4215);
CN_in_sig(542)	<=	VN_out_sig(4216);
CN_in_sig(2518)	<=	VN_out_sig(4217);
CN_in_sig(2918)	<=	VN_out_sig(4218);
CN_in_sig(4270)	<=	VN_out_sig(4219);
CN_in_sig(550)	<=	VN_out_sig(4220);
CN_in_sig(2526)	<=	VN_out_sig(4221);
CN_in_sig(2926)	<=	VN_out_sig(4222);
CN_in_sig(4278)	<=	VN_out_sig(4223);
CN_in_sig(558)	<=	VN_out_sig(4224);
CN_in_sig(2534)	<=	VN_out_sig(4225);
CN_in_sig(2934)	<=	VN_out_sig(4226);
CN_in_sig(4286)	<=	VN_out_sig(4227);
CN_in_sig(566)	<=	VN_out_sig(4228);
CN_in_sig(2542)	<=	VN_out_sig(4229);
CN_in_sig(2942)	<=	VN_out_sig(4230);
CN_in_sig(4294)	<=	VN_out_sig(4231);
CN_in_sig(574)	<=	VN_out_sig(4232);
CN_in_sig(2550)	<=	VN_out_sig(4233);
CN_in_sig(2950)	<=	VN_out_sig(4234);
CN_in_sig(4302)	<=	VN_out_sig(4235);
CN_in_sig(582)	<=	VN_out_sig(4236);
CN_in_sig(2558)	<=	VN_out_sig(4237);
CN_in_sig(2958)	<=	VN_out_sig(4238);
CN_in_sig(4310)	<=	VN_out_sig(4239);
CN_in_sig(590)	<=	VN_out_sig(4240);
CN_in_sig(2566)	<=	VN_out_sig(4241);
CN_in_sig(2966)	<=	VN_out_sig(4242);
CN_in_sig(4318)	<=	VN_out_sig(4243);
CN_in_sig(598)	<=	VN_out_sig(4244);
CN_in_sig(2574)	<=	VN_out_sig(4245);
CN_in_sig(2974)	<=	VN_out_sig(4246);
CN_in_sig(3894)	<=	VN_out_sig(4247);
CN_in_sig(606)	<=	VN_out_sig(4248);
CN_in_sig(2582)	<=	VN_out_sig(4249);
CN_in_sig(2982)	<=	VN_out_sig(4250);
CN_in_sig(3902)	<=	VN_out_sig(4251);
CN_in_sig(614)	<=	VN_out_sig(4252);
CN_in_sig(2590)	<=	VN_out_sig(4253);
CN_in_sig(2990)	<=	VN_out_sig(4254);
CN_in_sig(3910)	<=	VN_out_sig(4255);
CN_in_sig(622)	<=	VN_out_sig(4256);
CN_in_sig(2166)	<=	VN_out_sig(4257);
CN_in_sig(2998)	<=	VN_out_sig(4258);
CN_in_sig(3918)	<=	VN_out_sig(4259);
CN_in_sig(630)	<=	VN_out_sig(4260);
CN_in_sig(2174)	<=	VN_out_sig(4261);
CN_in_sig(3006)	<=	VN_out_sig(4262);
CN_in_sig(3926)	<=	VN_out_sig(4263);
CN_in_sig(638)	<=	VN_out_sig(4264);
CN_in_sig(2182)	<=	VN_out_sig(4265);
CN_in_sig(3014)	<=	VN_out_sig(4266);
CN_in_sig(3934)	<=	VN_out_sig(4267);
CN_in_sig(646)	<=	VN_out_sig(4268);
CN_in_sig(2190)	<=	VN_out_sig(4269);
CN_in_sig(3022)	<=	VN_out_sig(4270);
CN_in_sig(3942)	<=	VN_out_sig(4271);
CN_in_sig(654)	<=	VN_out_sig(4272);
CN_in_sig(2198)	<=	VN_out_sig(4273);
CN_in_sig(2598)	<=	VN_out_sig(4274);
CN_in_sig(3950)	<=	VN_out_sig(4275);
CN_in_sig(662)	<=	VN_out_sig(4276);
CN_in_sig(2206)	<=	VN_out_sig(4277);
CN_in_sig(2606)	<=	VN_out_sig(4278);
CN_in_sig(3958)	<=	VN_out_sig(4279);
CN_in_sig(670)	<=	VN_out_sig(4280);
CN_in_sig(2214)	<=	VN_out_sig(4281);
CN_in_sig(2614)	<=	VN_out_sig(4282);
CN_in_sig(3966)	<=	VN_out_sig(4283);
CN_in_sig(678)	<=	VN_out_sig(4284);
CN_in_sig(2222)	<=	VN_out_sig(4285);
CN_in_sig(2622)	<=	VN_out_sig(4286);
CN_in_sig(3974)	<=	VN_out_sig(4287);
CN_in_sig(686)	<=	VN_out_sig(4288);
CN_in_sig(2230)	<=	VN_out_sig(4289);
CN_in_sig(2630)	<=	VN_out_sig(4290);
CN_in_sig(3982)	<=	VN_out_sig(4291);
CN_in_sig(694)	<=	VN_out_sig(4292);
CN_in_sig(2238)	<=	VN_out_sig(4293);
CN_in_sig(2638)	<=	VN_out_sig(4294);
CN_in_sig(3990)	<=	VN_out_sig(4295);
CN_in_sig(702)	<=	VN_out_sig(4296);
CN_in_sig(2246)	<=	VN_out_sig(4297);
CN_in_sig(2646)	<=	VN_out_sig(4298);
CN_in_sig(3998)	<=	VN_out_sig(4299);
CN_in_sig(710)	<=	VN_out_sig(4300);
CN_in_sig(2254)	<=	VN_out_sig(4301);
CN_in_sig(2654)	<=	VN_out_sig(4302);
CN_in_sig(4006)	<=	VN_out_sig(4303);
CN_in_sig(718)	<=	VN_out_sig(4304);
CN_in_sig(2262)	<=	VN_out_sig(4305);
CN_in_sig(2662)	<=	VN_out_sig(4306);
CN_in_sig(4014)	<=	VN_out_sig(4307);
CN_in_sig(726)	<=	VN_out_sig(4308);
CN_in_sig(2270)	<=	VN_out_sig(4309);
CN_in_sig(2670)	<=	VN_out_sig(4310);
CN_in_sig(4022)	<=	VN_out_sig(4311);
CN_in_sig(734)	<=	VN_out_sig(4312);
CN_in_sig(2278)	<=	VN_out_sig(4313);
CN_in_sig(2678)	<=	VN_out_sig(4314);
CN_in_sig(4030)	<=	VN_out_sig(4315);
CN_in_sig(742)	<=	VN_out_sig(4316);
CN_in_sig(2286)	<=	VN_out_sig(4317);
CN_in_sig(2686)	<=	VN_out_sig(4318);
CN_in_sig(4038)	<=	VN_out_sig(4319);
CN_in_sig(1062)	<=	VN_out_sig(4320);
CN_in_sig(1806)	<=	VN_out_sig(4321);
CN_in_sig(3238)	<=	VN_out_sig(4322);
CN_in_sig(4470)	<=	VN_out_sig(4323);
CN_in_sig(1070)	<=	VN_out_sig(4324);
CN_in_sig(1814)	<=	VN_out_sig(4325);
CN_in_sig(3246)	<=	VN_out_sig(4326);
CN_in_sig(4478)	<=	VN_out_sig(4327);
CN_in_sig(1078)	<=	VN_out_sig(4328);
CN_in_sig(1822)	<=	VN_out_sig(4329);
CN_in_sig(3254)	<=	VN_out_sig(4330);
CN_in_sig(4486)	<=	VN_out_sig(4331);
CN_in_sig(1086)	<=	VN_out_sig(4332);
CN_in_sig(1830)	<=	VN_out_sig(4333);
CN_in_sig(3262)	<=	VN_out_sig(4334);
CN_in_sig(4494)	<=	VN_out_sig(4335);
CN_in_sig(1094)	<=	VN_out_sig(4336);
CN_in_sig(1838)	<=	VN_out_sig(4337);
CN_in_sig(3270)	<=	VN_out_sig(4338);
CN_in_sig(4502)	<=	VN_out_sig(4339);
CN_in_sig(1102)	<=	VN_out_sig(4340);
CN_in_sig(1846)	<=	VN_out_sig(4341);
CN_in_sig(3278)	<=	VN_out_sig(4342);
CN_in_sig(4510)	<=	VN_out_sig(4343);
CN_in_sig(1110)	<=	VN_out_sig(4344);
CN_in_sig(1854)	<=	VN_out_sig(4345);
CN_in_sig(3286)	<=	VN_out_sig(4346);
CN_in_sig(4518)	<=	VN_out_sig(4347);
CN_in_sig(1118)	<=	VN_out_sig(4348);
CN_in_sig(1862)	<=	VN_out_sig(4349);
CN_in_sig(3294)	<=	VN_out_sig(4350);
CN_in_sig(4526)	<=	VN_out_sig(4351);
CN_in_sig(1126)	<=	VN_out_sig(4352);
CN_in_sig(1870)	<=	VN_out_sig(4353);
CN_in_sig(3302)	<=	VN_out_sig(4354);
CN_in_sig(4534)	<=	VN_out_sig(4355);
CN_in_sig(1134)	<=	VN_out_sig(4356);
CN_in_sig(1878)	<=	VN_out_sig(4357);
CN_in_sig(3310)	<=	VN_out_sig(4358);
CN_in_sig(4542)	<=	VN_out_sig(4359);
CN_in_sig(1142)	<=	VN_out_sig(4360);
CN_in_sig(1886)	<=	VN_out_sig(4361);
CN_in_sig(3318)	<=	VN_out_sig(4362);
CN_in_sig(4550)	<=	VN_out_sig(4363);
CN_in_sig(1150)	<=	VN_out_sig(4364);
CN_in_sig(1894)	<=	VN_out_sig(4365);
CN_in_sig(3326)	<=	VN_out_sig(4366);
CN_in_sig(4558)	<=	VN_out_sig(4367);
CN_in_sig(1158)	<=	VN_out_sig(4368);
CN_in_sig(1902)	<=	VN_out_sig(4369);
CN_in_sig(3334)	<=	VN_out_sig(4370);
CN_in_sig(4566)	<=	VN_out_sig(4371);
CN_in_sig(1166)	<=	VN_out_sig(4372);
CN_in_sig(1910)	<=	VN_out_sig(4373);
CN_in_sig(3342)	<=	VN_out_sig(4374);
CN_in_sig(4574)	<=	VN_out_sig(4375);
CN_in_sig(1174)	<=	VN_out_sig(4376);
CN_in_sig(1918)	<=	VN_out_sig(4377);
CN_in_sig(3350)	<=	VN_out_sig(4378);
CN_in_sig(4582)	<=	VN_out_sig(4379);
CN_in_sig(1182)	<=	VN_out_sig(4380);
CN_in_sig(1926)	<=	VN_out_sig(4381);
CN_in_sig(3358)	<=	VN_out_sig(4382);
CN_in_sig(4590)	<=	VN_out_sig(4383);
CN_in_sig(1190)	<=	VN_out_sig(4384);
CN_in_sig(1934)	<=	VN_out_sig(4385);
CN_in_sig(3366)	<=	VN_out_sig(4386);
CN_in_sig(4598)	<=	VN_out_sig(4387);
CN_in_sig(1198)	<=	VN_out_sig(4388);
CN_in_sig(1942)	<=	VN_out_sig(4389);
CN_in_sig(3374)	<=	VN_out_sig(4390);
CN_in_sig(4606)	<=	VN_out_sig(4391);
CN_in_sig(1206)	<=	VN_out_sig(4392);
CN_in_sig(1950)	<=	VN_out_sig(4393);
CN_in_sig(3382)	<=	VN_out_sig(4394);
CN_in_sig(4614)	<=	VN_out_sig(4395);
CN_in_sig(1214)	<=	VN_out_sig(4396);
CN_in_sig(1958)	<=	VN_out_sig(4397);
CN_in_sig(3390)	<=	VN_out_sig(4398);
CN_in_sig(4622)	<=	VN_out_sig(4399);
CN_in_sig(1222)	<=	VN_out_sig(4400);
CN_in_sig(1966)	<=	VN_out_sig(4401);
CN_in_sig(3398)	<=	VN_out_sig(4402);
CN_in_sig(4630)	<=	VN_out_sig(4403);
CN_in_sig(1230)	<=	VN_out_sig(4404);
CN_in_sig(1974)	<=	VN_out_sig(4405);
CN_in_sig(3406)	<=	VN_out_sig(4406);
CN_in_sig(4638)	<=	VN_out_sig(4407);
CN_in_sig(1238)	<=	VN_out_sig(4408);
CN_in_sig(1982)	<=	VN_out_sig(4409);
CN_in_sig(3414)	<=	VN_out_sig(4410);
CN_in_sig(4646)	<=	VN_out_sig(4411);
CN_in_sig(1246)	<=	VN_out_sig(4412);
CN_in_sig(1990)	<=	VN_out_sig(4413);
CN_in_sig(3422)	<=	VN_out_sig(4414);
CN_in_sig(4654)	<=	VN_out_sig(4415);
CN_in_sig(1254)	<=	VN_out_sig(4416);
CN_in_sig(1998)	<=	VN_out_sig(4417);
CN_in_sig(3430)	<=	VN_out_sig(4418);
CN_in_sig(4662)	<=	VN_out_sig(4419);
CN_in_sig(1262)	<=	VN_out_sig(4420);
CN_in_sig(2006)	<=	VN_out_sig(4421);
CN_in_sig(3438)	<=	VN_out_sig(4422);
CN_in_sig(4670)	<=	VN_out_sig(4423);
CN_in_sig(1270)	<=	VN_out_sig(4424);
CN_in_sig(2014)	<=	VN_out_sig(4425);
CN_in_sig(3446)	<=	VN_out_sig(4426);
CN_in_sig(4678)	<=	VN_out_sig(4427);
CN_in_sig(1278)	<=	VN_out_sig(4428);
CN_in_sig(2022)	<=	VN_out_sig(4429);
CN_in_sig(3454)	<=	VN_out_sig(4430);
CN_in_sig(4686)	<=	VN_out_sig(4431);
CN_in_sig(1286)	<=	VN_out_sig(4432);
CN_in_sig(2030)	<=	VN_out_sig(4433);
CN_in_sig(3030)	<=	VN_out_sig(4434);
CN_in_sig(4694)	<=	VN_out_sig(4435);
CN_in_sig(1294)	<=	VN_out_sig(4436);
CN_in_sig(2038)	<=	VN_out_sig(4437);
CN_in_sig(3038)	<=	VN_out_sig(4438);
CN_in_sig(4702)	<=	VN_out_sig(4439);
CN_in_sig(870)	<=	VN_out_sig(4440);
CN_in_sig(2046)	<=	VN_out_sig(4441);
CN_in_sig(3046)	<=	VN_out_sig(4442);
CN_in_sig(4710)	<=	VN_out_sig(4443);
CN_in_sig(878)	<=	VN_out_sig(4444);
CN_in_sig(2054)	<=	VN_out_sig(4445);
CN_in_sig(3054)	<=	VN_out_sig(4446);
CN_in_sig(4718)	<=	VN_out_sig(4447);
CN_in_sig(886)	<=	VN_out_sig(4448);
CN_in_sig(2062)	<=	VN_out_sig(4449);
CN_in_sig(3062)	<=	VN_out_sig(4450);
CN_in_sig(4726)	<=	VN_out_sig(4451);
CN_in_sig(894)	<=	VN_out_sig(4452);
CN_in_sig(2070)	<=	VN_out_sig(4453);
CN_in_sig(3070)	<=	VN_out_sig(4454);
CN_in_sig(4734)	<=	VN_out_sig(4455);
CN_in_sig(902)	<=	VN_out_sig(4456);
CN_in_sig(2078)	<=	VN_out_sig(4457);
CN_in_sig(3078)	<=	VN_out_sig(4458);
CN_in_sig(4742)	<=	VN_out_sig(4459);
CN_in_sig(910)	<=	VN_out_sig(4460);
CN_in_sig(2086)	<=	VN_out_sig(4461);
CN_in_sig(3086)	<=	VN_out_sig(4462);
CN_in_sig(4750)	<=	VN_out_sig(4463);
CN_in_sig(918)	<=	VN_out_sig(4464);
CN_in_sig(2094)	<=	VN_out_sig(4465);
CN_in_sig(3094)	<=	VN_out_sig(4466);
CN_in_sig(4326)	<=	VN_out_sig(4467);
CN_in_sig(926)	<=	VN_out_sig(4468);
CN_in_sig(2102)	<=	VN_out_sig(4469);
CN_in_sig(3102)	<=	VN_out_sig(4470);
CN_in_sig(4334)	<=	VN_out_sig(4471);
CN_in_sig(934)	<=	VN_out_sig(4472);
CN_in_sig(2110)	<=	VN_out_sig(4473);
CN_in_sig(3110)	<=	VN_out_sig(4474);
CN_in_sig(4342)	<=	VN_out_sig(4475);
CN_in_sig(942)	<=	VN_out_sig(4476);
CN_in_sig(2118)	<=	VN_out_sig(4477);
CN_in_sig(3118)	<=	VN_out_sig(4478);
CN_in_sig(4350)	<=	VN_out_sig(4479);
CN_in_sig(950)	<=	VN_out_sig(4480);
CN_in_sig(2126)	<=	VN_out_sig(4481);
CN_in_sig(3126)	<=	VN_out_sig(4482);
CN_in_sig(4358)	<=	VN_out_sig(4483);
CN_in_sig(958)	<=	VN_out_sig(4484);
CN_in_sig(2134)	<=	VN_out_sig(4485);
CN_in_sig(3134)	<=	VN_out_sig(4486);
CN_in_sig(4366)	<=	VN_out_sig(4487);
CN_in_sig(966)	<=	VN_out_sig(4488);
CN_in_sig(2142)	<=	VN_out_sig(4489);
CN_in_sig(3142)	<=	VN_out_sig(4490);
CN_in_sig(4374)	<=	VN_out_sig(4491);
CN_in_sig(974)	<=	VN_out_sig(4492);
CN_in_sig(2150)	<=	VN_out_sig(4493);
CN_in_sig(3150)	<=	VN_out_sig(4494);
CN_in_sig(4382)	<=	VN_out_sig(4495);
CN_in_sig(982)	<=	VN_out_sig(4496);
CN_in_sig(2158)	<=	VN_out_sig(4497);
CN_in_sig(3158)	<=	VN_out_sig(4498);
CN_in_sig(4390)	<=	VN_out_sig(4499);
CN_in_sig(990)	<=	VN_out_sig(4500);
CN_in_sig(1734)	<=	VN_out_sig(4501);
CN_in_sig(3166)	<=	VN_out_sig(4502);
CN_in_sig(4398)	<=	VN_out_sig(4503);
CN_in_sig(998)	<=	VN_out_sig(4504);
CN_in_sig(1742)	<=	VN_out_sig(4505);
CN_in_sig(3174)	<=	VN_out_sig(4506);
CN_in_sig(4406)	<=	VN_out_sig(4507);
CN_in_sig(1006)	<=	VN_out_sig(4508);
CN_in_sig(1750)	<=	VN_out_sig(4509);
CN_in_sig(3182)	<=	VN_out_sig(4510);
CN_in_sig(4414)	<=	VN_out_sig(4511);
CN_in_sig(1014)	<=	VN_out_sig(4512);
CN_in_sig(1758)	<=	VN_out_sig(4513);
CN_in_sig(3190)	<=	VN_out_sig(4514);
CN_in_sig(4422)	<=	VN_out_sig(4515);
CN_in_sig(1022)	<=	VN_out_sig(4516);
CN_in_sig(1766)	<=	VN_out_sig(4517);
CN_in_sig(3198)	<=	VN_out_sig(4518);
CN_in_sig(4430)	<=	VN_out_sig(4519);
CN_in_sig(1030)	<=	VN_out_sig(4520);
CN_in_sig(1774)	<=	VN_out_sig(4521);
CN_in_sig(3206)	<=	VN_out_sig(4522);
CN_in_sig(4438)	<=	VN_out_sig(4523);
CN_in_sig(1038)	<=	VN_out_sig(4524);
CN_in_sig(1782)	<=	VN_out_sig(4525);
CN_in_sig(3214)	<=	VN_out_sig(4526);
CN_in_sig(4446)	<=	VN_out_sig(4527);
CN_in_sig(1046)	<=	VN_out_sig(4528);
CN_in_sig(1790)	<=	VN_out_sig(4529);
CN_in_sig(3222)	<=	VN_out_sig(4530);
CN_in_sig(4454)	<=	VN_out_sig(4531);
CN_in_sig(1054)	<=	VN_out_sig(4532);
CN_in_sig(1798)	<=	VN_out_sig(4533);
CN_in_sig(3230)	<=	VN_out_sig(4534);
CN_in_sig(4462)	<=	VN_out_sig(4535);
CN_in_sig(1039)	<=	VN_out_sig(4536);
CN_in_sig(2031)	<=	VN_out_sig(4537);
CN_in_sig(3135)	<=	VN_out_sig(4538);
CN_in_sig(4455)	<=	VN_out_sig(4539);
CN_in_sig(1047)	<=	VN_out_sig(4540);
CN_in_sig(2039)	<=	VN_out_sig(4541);
CN_in_sig(3143)	<=	VN_out_sig(4542);
CN_in_sig(4463)	<=	VN_out_sig(4543);
CN_in_sig(1055)	<=	VN_out_sig(4544);
CN_in_sig(2047)	<=	VN_out_sig(4545);
CN_in_sig(3151)	<=	VN_out_sig(4546);
CN_in_sig(4471)	<=	VN_out_sig(4547);
CN_in_sig(1063)	<=	VN_out_sig(4548);
CN_in_sig(2055)	<=	VN_out_sig(4549);
CN_in_sig(3159)	<=	VN_out_sig(4550);
CN_in_sig(4479)	<=	VN_out_sig(4551);
CN_in_sig(1071)	<=	VN_out_sig(4552);
CN_in_sig(2063)	<=	VN_out_sig(4553);
CN_in_sig(3167)	<=	VN_out_sig(4554);
CN_in_sig(4487)	<=	VN_out_sig(4555);
CN_in_sig(1079)	<=	VN_out_sig(4556);
CN_in_sig(2071)	<=	VN_out_sig(4557);
CN_in_sig(3175)	<=	VN_out_sig(4558);
CN_in_sig(4495)	<=	VN_out_sig(4559);
CN_in_sig(1087)	<=	VN_out_sig(4560);
CN_in_sig(2079)	<=	VN_out_sig(4561);
CN_in_sig(3183)	<=	VN_out_sig(4562);
CN_in_sig(4503)	<=	VN_out_sig(4563);
CN_in_sig(1095)	<=	VN_out_sig(4564);
CN_in_sig(2087)	<=	VN_out_sig(4565);
CN_in_sig(3191)	<=	VN_out_sig(4566);
CN_in_sig(4511)	<=	VN_out_sig(4567);
CN_in_sig(1103)	<=	VN_out_sig(4568);
CN_in_sig(2095)	<=	VN_out_sig(4569);
CN_in_sig(3199)	<=	VN_out_sig(4570);
CN_in_sig(4519)	<=	VN_out_sig(4571);
CN_in_sig(1111)	<=	VN_out_sig(4572);
CN_in_sig(2103)	<=	VN_out_sig(4573);
CN_in_sig(3207)	<=	VN_out_sig(4574);
CN_in_sig(4527)	<=	VN_out_sig(4575);
CN_in_sig(1119)	<=	VN_out_sig(4576);
CN_in_sig(2111)	<=	VN_out_sig(4577);
CN_in_sig(3215)	<=	VN_out_sig(4578);
CN_in_sig(4535)	<=	VN_out_sig(4579);
CN_in_sig(1127)	<=	VN_out_sig(4580);
CN_in_sig(2119)	<=	VN_out_sig(4581);
CN_in_sig(3223)	<=	VN_out_sig(4582);
CN_in_sig(4543)	<=	VN_out_sig(4583);
CN_in_sig(1135)	<=	VN_out_sig(4584);
CN_in_sig(2127)	<=	VN_out_sig(4585);
CN_in_sig(3231)	<=	VN_out_sig(4586);
CN_in_sig(4551)	<=	VN_out_sig(4587);
CN_in_sig(1143)	<=	VN_out_sig(4588);
CN_in_sig(2135)	<=	VN_out_sig(4589);
CN_in_sig(3239)	<=	VN_out_sig(4590);
CN_in_sig(4559)	<=	VN_out_sig(4591);
CN_in_sig(1151)	<=	VN_out_sig(4592);
CN_in_sig(2143)	<=	VN_out_sig(4593);
CN_in_sig(3247)	<=	VN_out_sig(4594);
CN_in_sig(4567)	<=	VN_out_sig(4595);
CN_in_sig(1159)	<=	VN_out_sig(4596);
CN_in_sig(2151)	<=	VN_out_sig(4597);
CN_in_sig(3255)	<=	VN_out_sig(4598);
CN_in_sig(4575)	<=	VN_out_sig(4599);
CN_in_sig(1167)	<=	VN_out_sig(4600);
CN_in_sig(2159)	<=	VN_out_sig(4601);
CN_in_sig(3263)	<=	VN_out_sig(4602);
CN_in_sig(4583)	<=	VN_out_sig(4603);
CN_in_sig(1175)	<=	VN_out_sig(4604);
CN_in_sig(1735)	<=	VN_out_sig(4605);
CN_in_sig(3271)	<=	VN_out_sig(4606);
CN_in_sig(4591)	<=	VN_out_sig(4607);
CN_in_sig(1183)	<=	VN_out_sig(4608);
CN_in_sig(1743)	<=	VN_out_sig(4609);
CN_in_sig(3279)	<=	VN_out_sig(4610);
CN_in_sig(4599)	<=	VN_out_sig(4611);
CN_in_sig(1191)	<=	VN_out_sig(4612);
CN_in_sig(1751)	<=	VN_out_sig(4613);
CN_in_sig(3287)	<=	VN_out_sig(4614);
CN_in_sig(4607)	<=	VN_out_sig(4615);
CN_in_sig(1199)	<=	VN_out_sig(4616);
CN_in_sig(1759)	<=	VN_out_sig(4617);
CN_in_sig(3295)	<=	VN_out_sig(4618);
CN_in_sig(4615)	<=	VN_out_sig(4619);
CN_in_sig(1207)	<=	VN_out_sig(4620);
CN_in_sig(1767)	<=	VN_out_sig(4621);
CN_in_sig(3303)	<=	VN_out_sig(4622);
CN_in_sig(4623)	<=	VN_out_sig(4623);
CN_in_sig(1215)	<=	VN_out_sig(4624);
CN_in_sig(1775)	<=	VN_out_sig(4625);
CN_in_sig(3311)	<=	VN_out_sig(4626);
CN_in_sig(4631)	<=	VN_out_sig(4627);
CN_in_sig(1223)	<=	VN_out_sig(4628);
CN_in_sig(1783)	<=	VN_out_sig(4629);
CN_in_sig(3319)	<=	VN_out_sig(4630);
CN_in_sig(4639)	<=	VN_out_sig(4631);
CN_in_sig(1231)	<=	VN_out_sig(4632);
CN_in_sig(1791)	<=	VN_out_sig(4633);
CN_in_sig(3327)	<=	VN_out_sig(4634);
CN_in_sig(4647)	<=	VN_out_sig(4635);
CN_in_sig(1239)	<=	VN_out_sig(4636);
CN_in_sig(1799)	<=	VN_out_sig(4637);
CN_in_sig(3335)	<=	VN_out_sig(4638);
CN_in_sig(4655)	<=	VN_out_sig(4639);
CN_in_sig(1247)	<=	VN_out_sig(4640);
CN_in_sig(1807)	<=	VN_out_sig(4641);
CN_in_sig(3343)	<=	VN_out_sig(4642);
CN_in_sig(4663)	<=	VN_out_sig(4643);
CN_in_sig(1255)	<=	VN_out_sig(4644);
CN_in_sig(1815)	<=	VN_out_sig(4645);
CN_in_sig(3351)	<=	VN_out_sig(4646);
CN_in_sig(4671)	<=	VN_out_sig(4647);
CN_in_sig(1263)	<=	VN_out_sig(4648);
CN_in_sig(1823)	<=	VN_out_sig(4649);
CN_in_sig(3359)	<=	VN_out_sig(4650);
CN_in_sig(4679)	<=	VN_out_sig(4651);
CN_in_sig(1271)	<=	VN_out_sig(4652);
CN_in_sig(1831)	<=	VN_out_sig(4653);
CN_in_sig(3367)	<=	VN_out_sig(4654);
CN_in_sig(4687)	<=	VN_out_sig(4655);
CN_in_sig(1279)	<=	VN_out_sig(4656);
CN_in_sig(1839)	<=	VN_out_sig(4657);
CN_in_sig(3375)	<=	VN_out_sig(4658);
CN_in_sig(4695)	<=	VN_out_sig(4659);
CN_in_sig(1287)	<=	VN_out_sig(4660);
CN_in_sig(1847)	<=	VN_out_sig(4661);
CN_in_sig(3383)	<=	VN_out_sig(4662);
CN_in_sig(4703)	<=	VN_out_sig(4663);
CN_in_sig(1295)	<=	VN_out_sig(4664);
CN_in_sig(1855)	<=	VN_out_sig(4665);
CN_in_sig(3391)	<=	VN_out_sig(4666);
CN_in_sig(4711)	<=	VN_out_sig(4667);
CN_in_sig(871)	<=	VN_out_sig(4668);
CN_in_sig(1863)	<=	VN_out_sig(4669);
CN_in_sig(3399)	<=	VN_out_sig(4670);
CN_in_sig(4719)	<=	VN_out_sig(4671);
CN_in_sig(879)	<=	VN_out_sig(4672);
CN_in_sig(1871)	<=	VN_out_sig(4673);
CN_in_sig(3407)	<=	VN_out_sig(4674);
CN_in_sig(4727)	<=	VN_out_sig(4675);
CN_in_sig(887)	<=	VN_out_sig(4676);
CN_in_sig(1879)	<=	VN_out_sig(4677);
CN_in_sig(3415)	<=	VN_out_sig(4678);
CN_in_sig(4735)	<=	VN_out_sig(4679);
CN_in_sig(895)	<=	VN_out_sig(4680);
CN_in_sig(1887)	<=	VN_out_sig(4681);
CN_in_sig(3423)	<=	VN_out_sig(4682);
CN_in_sig(4743)	<=	VN_out_sig(4683);
CN_in_sig(903)	<=	VN_out_sig(4684);
CN_in_sig(1895)	<=	VN_out_sig(4685);
CN_in_sig(3431)	<=	VN_out_sig(4686);
CN_in_sig(4751)	<=	VN_out_sig(4687);
CN_in_sig(911)	<=	VN_out_sig(4688);
CN_in_sig(1903)	<=	VN_out_sig(4689);
CN_in_sig(3439)	<=	VN_out_sig(4690);
CN_in_sig(4327)	<=	VN_out_sig(4691);
CN_in_sig(919)	<=	VN_out_sig(4692);
CN_in_sig(1911)	<=	VN_out_sig(4693);
CN_in_sig(3447)	<=	VN_out_sig(4694);
CN_in_sig(4335)	<=	VN_out_sig(4695);
CN_in_sig(927)	<=	VN_out_sig(4696);
CN_in_sig(1919)	<=	VN_out_sig(4697);
CN_in_sig(3455)	<=	VN_out_sig(4698);
CN_in_sig(4343)	<=	VN_out_sig(4699);
CN_in_sig(935)	<=	VN_out_sig(4700);
CN_in_sig(1927)	<=	VN_out_sig(4701);
CN_in_sig(3031)	<=	VN_out_sig(4702);
CN_in_sig(4351)	<=	VN_out_sig(4703);
CN_in_sig(943)	<=	VN_out_sig(4704);
CN_in_sig(1935)	<=	VN_out_sig(4705);
CN_in_sig(3039)	<=	VN_out_sig(4706);
CN_in_sig(4359)	<=	VN_out_sig(4707);
CN_in_sig(951)	<=	VN_out_sig(4708);
CN_in_sig(1943)	<=	VN_out_sig(4709);
CN_in_sig(3047)	<=	VN_out_sig(4710);
CN_in_sig(4367)	<=	VN_out_sig(4711);
CN_in_sig(959)	<=	VN_out_sig(4712);
CN_in_sig(1951)	<=	VN_out_sig(4713);
CN_in_sig(3055)	<=	VN_out_sig(4714);
CN_in_sig(4375)	<=	VN_out_sig(4715);
CN_in_sig(967)	<=	VN_out_sig(4716);
CN_in_sig(1959)	<=	VN_out_sig(4717);
CN_in_sig(3063)	<=	VN_out_sig(4718);
CN_in_sig(4383)	<=	VN_out_sig(4719);
CN_in_sig(975)	<=	VN_out_sig(4720);
CN_in_sig(1967)	<=	VN_out_sig(4721);
CN_in_sig(3071)	<=	VN_out_sig(4722);
CN_in_sig(4391)	<=	VN_out_sig(4723);
CN_in_sig(983)	<=	VN_out_sig(4724);
CN_in_sig(1975)	<=	VN_out_sig(4725);
CN_in_sig(3079)	<=	VN_out_sig(4726);
CN_in_sig(4399)	<=	VN_out_sig(4727);
CN_in_sig(991)	<=	VN_out_sig(4728);
CN_in_sig(1983)	<=	VN_out_sig(4729);
CN_in_sig(3087)	<=	VN_out_sig(4730);
CN_in_sig(4407)	<=	VN_out_sig(4731);
CN_in_sig(999)	<=	VN_out_sig(4732);
CN_in_sig(1991)	<=	VN_out_sig(4733);
CN_in_sig(3095)	<=	VN_out_sig(4734);
CN_in_sig(4415)	<=	VN_out_sig(4735);
CN_in_sig(1007)	<=	VN_out_sig(4736);
CN_in_sig(1999)	<=	VN_out_sig(4737);
CN_in_sig(3103)	<=	VN_out_sig(4738);
CN_in_sig(4423)	<=	VN_out_sig(4739);
CN_in_sig(1015)	<=	VN_out_sig(4740);
CN_in_sig(2007)	<=	VN_out_sig(4741);
CN_in_sig(3111)	<=	VN_out_sig(4742);
CN_in_sig(4431)	<=	VN_out_sig(4743);
CN_in_sig(1023)	<=	VN_out_sig(4744);
CN_in_sig(2015)	<=	VN_out_sig(4745);
CN_in_sig(3119)	<=	VN_out_sig(4746);
CN_in_sig(4439)	<=	VN_out_sig(4747);
CN_in_sig(1031)	<=	VN_out_sig(4748);
CN_in_sig(2023)	<=	VN_out_sig(4749);
CN_in_sig(3127)	<=	VN_out_sig(4750);
CN_in_sig(4447)	<=	VN_out_sig(4751);
CN_in_sig(735)	<=	VN_out_sig(4752);
CN_in_sig(2351)	<=	VN_out_sig(4753);
CN_in_sig(2719)	<=	VN_out_sig(4754);
CN_in_sig(3975)	<=	VN_out_sig(4755);
CN_in_sig(743)	<=	VN_out_sig(4756);
CN_in_sig(2359)	<=	VN_out_sig(4757);
CN_in_sig(2727)	<=	VN_out_sig(4758);
CN_in_sig(3983)	<=	VN_out_sig(4759);
CN_in_sig(751)	<=	VN_out_sig(4760);
CN_in_sig(2367)	<=	VN_out_sig(4761);
CN_in_sig(2735)	<=	VN_out_sig(4762);
CN_in_sig(3991)	<=	VN_out_sig(4763);
CN_in_sig(759)	<=	VN_out_sig(4764);
CN_in_sig(2375)	<=	VN_out_sig(4765);
CN_in_sig(2743)	<=	VN_out_sig(4766);
CN_in_sig(3999)	<=	VN_out_sig(4767);
CN_in_sig(767)	<=	VN_out_sig(4768);
CN_in_sig(2383)	<=	VN_out_sig(4769);
CN_in_sig(2751)	<=	VN_out_sig(4770);
CN_in_sig(4007)	<=	VN_out_sig(4771);
CN_in_sig(775)	<=	VN_out_sig(4772);
CN_in_sig(2391)	<=	VN_out_sig(4773);
CN_in_sig(2759)	<=	VN_out_sig(4774);
CN_in_sig(4015)	<=	VN_out_sig(4775);
CN_in_sig(783)	<=	VN_out_sig(4776);
CN_in_sig(2399)	<=	VN_out_sig(4777);
CN_in_sig(2767)	<=	VN_out_sig(4778);
CN_in_sig(4023)	<=	VN_out_sig(4779);
CN_in_sig(791)	<=	VN_out_sig(4780);
CN_in_sig(2407)	<=	VN_out_sig(4781);
CN_in_sig(2775)	<=	VN_out_sig(4782);
CN_in_sig(4031)	<=	VN_out_sig(4783);
CN_in_sig(799)	<=	VN_out_sig(4784);
CN_in_sig(2415)	<=	VN_out_sig(4785);
CN_in_sig(2783)	<=	VN_out_sig(4786);
CN_in_sig(4039)	<=	VN_out_sig(4787);
CN_in_sig(807)	<=	VN_out_sig(4788);
CN_in_sig(2423)	<=	VN_out_sig(4789);
CN_in_sig(2791)	<=	VN_out_sig(4790);
CN_in_sig(4047)	<=	VN_out_sig(4791);
CN_in_sig(815)	<=	VN_out_sig(4792);
CN_in_sig(2431)	<=	VN_out_sig(4793);
CN_in_sig(2799)	<=	VN_out_sig(4794);
CN_in_sig(4055)	<=	VN_out_sig(4795);
CN_in_sig(823)	<=	VN_out_sig(4796);
CN_in_sig(2439)	<=	VN_out_sig(4797);
CN_in_sig(2807)	<=	VN_out_sig(4798);
CN_in_sig(4063)	<=	VN_out_sig(4799);
CN_in_sig(831)	<=	VN_out_sig(4800);
CN_in_sig(2447)	<=	VN_out_sig(4801);
CN_in_sig(2815)	<=	VN_out_sig(4802);
CN_in_sig(4071)	<=	VN_out_sig(4803);
CN_in_sig(839)	<=	VN_out_sig(4804);
CN_in_sig(2455)	<=	VN_out_sig(4805);
CN_in_sig(2823)	<=	VN_out_sig(4806);
CN_in_sig(4079)	<=	VN_out_sig(4807);
CN_in_sig(847)	<=	VN_out_sig(4808);
CN_in_sig(2463)	<=	VN_out_sig(4809);
CN_in_sig(2831)	<=	VN_out_sig(4810);
CN_in_sig(4087)	<=	VN_out_sig(4811);
CN_in_sig(855)	<=	VN_out_sig(4812);
CN_in_sig(2471)	<=	VN_out_sig(4813);
CN_in_sig(2839)	<=	VN_out_sig(4814);
CN_in_sig(4095)	<=	VN_out_sig(4815);
CN_in_sig(863)	<=	VN_out_sig(4816);
CN_in_sig(2479)	<=	VN_out_sig(4817);
CN_in_sig(2847)	<=	VN_out_sig(4818);
CN_in_sig(4103)	<=	VN_out_sig(4819);
CN_in_sig(439)	<=	VN_out_sig(4820);
CN_in_sig(2487)	<=	VN_out_sig(4821);
CN_in_sig(2855)	<=	VN_out_sig(4822);
CN_in_sig(4111)	<=	VN_out_sig(4823);
CN_in_sig(447)	<=	VN_out_sig(4824);
CN_in_sig(2495)	<=	VN_out_sig(4825);
CN_in_sig(2863)	<=	VN_out_sig(4826);
CN_in_sig(4119)	<=	VN_out_sig(4827);
CN_in_sig(455)	<=	VN_out_sig(4828);
CN_in_sig(2503)	<=	VN_out_sig(4829);
CN_in_sig(2871)	<=	VN_out_sig(4830);
CN_in_sig(4127)	<=	VN_out_sig(4831);
CN_in_sig(463)	<=	VN_out_sig(4832);
CN_in_sig(2511)	<=	VN_out_sig(4833);
CN_in_sig(2879)	<=	VN_out_sig(4834);
CN_in_sig(4135)	<=	VN_out_sig(4835);
CN_in_sig(471)	<=	VN_out_sig(4836);
CN_in_sig(2519)	<=	VN_out_sig(4837);
CN_in_sig(2887)	<=	VN_out_sig(4838);
CN_in_sig(4143)	<=	VN_out_sig(4839);
CN_in_sig(479)	<=	VN_out_sig(4840);
CN_in_sig(2527)	<=	VN_out_sig(4841);
CN_in_sig(2895)	<=	VN_out_sig(4842);
CN_in_sig(4151)	<=	VN_out_sig(4843);
CN_in_sig(487)	<=	VN_out_sig(4844);
CN_in_sig(2535)	<=	VN_out_sig(4845);
CN_in_sig(2903)	<=	VN_out_sig(4846);
CN_in_sig(4159)	<=	VN_out_sig(4847);
CN_in_sig(495)	<=	VN_out_sig(4848);
CN_in_sig(2543)	<=	VN_out_sig(4849);
CN_in_sig(2911)	<=	VN_out_sig(4850);
CN_in_sig(4167)	<=	VN_out_sig(4851);
CN_in_sig(503)	<=	VN_out_sig(4852);
CN_in_sig(2551)	<=	VN_out_sig(4853);
CN_in_sig(2919)	<=	VN_out_sig(4854);
CN_in_sig(4175)	<=	VN_out_sig(4855);
CN_in_sig(511)	<=	VN_out_sig(4856);
CN_in_sig(2559)	<=	VN_out_sig(4857);
CN_in_sig(2927)	<=	VN_out_sig(4858);
CN_in_sig(4183)	<=	VN_out_sig(4859);
CN_in_sig(519)	<=	VN_out_sig(4860);
CN_in_sig(2567)	<=	VN_out_sig(4861);
CN_in_sig(2935)	<=	VN_out_sig(4862);
CN_in_sig(4191)	<=	VN_out_sig(4863);
CN_in_sig(527)	<=	VN_out_sig(4864);
CN_in_sig(2575)	<=	VN_out_sig(4865);
CN_in_sig(2943)	<=	VN_out_sig(4866);
CN_in_sig(4199)	<=	VN_out_sig(4867);
CN_in_sig(535)	<=	VN_out_sig(4868);
CN_in_sig(2583)	<=	VN_out_sig(4869);
CN_in_sig(2951)	<=	VN_out_sig(4870);
CN_in_sig(4207)	<=	VN_out_sig(4871);
CN_in_sig(543)	<=	VN_out_sig(4872);
CN_in_sig(2591)	<=	VN_out_sig(4873);
CN_in_sig(2959)	<=	VN_out_sig(4874);
CN_in_sig(4215)	<=	VN_out_sig(4875);
CN_in_sig(551)	<=	VN_out_sig(4876);
CN_in_sig(2167)	<=	VN_out_sig(4877);
CN_in_sig(2967)	<=	VN_out_sig(4878);
CN_in_sig(4223)	<=	VN_out_sig(4879);
CN_in_sig(559)	<=	VN_out_sig(4880);
CN_in_sig(2175)	<=	VN_out_sig(4881);
CN_in_sig(2975)	<=	VN_out_sig(4882);
CN_in_sig(4231)	<=	VN_out_sig(4883);
CN_in_sig(567)	<=	VN_out_sig(4884);
CN_in_sig(2183)	<=	VN_out_sig(4885);
CN_in_sig(2983)	<=	VN_out_sig(4886);
CN_in_sig(4239)	<=	VN_out_sig(4887);
CN_in_sig(575)	<=	VN_out_sig(4888);
CN_in_sig(2191)	<=	VN_out_sig(4889);
CN_in_sig(2991)	<=	VN_out_sig(4890);
CN_in_sig(4247)	<=	VN_out_sig(4891);
CN_in_sig(583)	<=	VN_out_sig(4892);
CN_in_sig(2199)	<=	VN_out_sig(4893);
CN_in_sig(2999)	<=	VN_out_sig(4894);
CN_in_sig(4255)	<=	VN_out_sig(4895);
CN_in_sig(591)	<=	VN_out_sig(4896);
CN_in_sig(2207)	<=	VN_out_sig(4897);
CN_in_sig(3007)	<=	VN_out_sig(4898);
CN_in_sig(4263)	<=	VN_out_sig(4899);
CN_in_sig(599)	<=	VN_out_sig(4900);
CN_in_sig(2215)	<=	VN_out_sig(4901);
CN_in_sig(3015)	<=	VN_out_sig(4902);
CN_in_sig(4271)	<=	VN_out_sig(4903);
CN_in_sig(607)	<=	VN_out_sig(4904);
CN_in_sig(2223)	<=	VN_out_sig(4905);
CN_in_sig(3023)	<=	VN_out_sig(4906);
CN_in_sig(4279)	<=	VN_out_sig(4907);
CN_in_sig(615)	<=	VN_out_sig(4908);
CN_in_sig(2231)	<=	VN_out_sig(4909);
CN_in_sig(2599)	<=	VN_out_sig(4910);
CN_in_sig(4287)	<=	VN_out_sig(4911);
CN_in_sig(623)	<=	VN_out_sig(4912);
CN_in_sig(2239)	<=	VN_out_sig(4913);
CN_in_sig(2607)	<=	VN_out_sig(4914);
CN_in_sig(4295)	<=	VN_out_sig(4915);
CN_in_sig(631)	<=	VN_out_sig(4916);
CN_in_sig(2247)	<=	VN_out_sig(4917);
CN_in_sig(2615)	<=	VN_out_sig(4918);
CN_in_sig(4303)	<=	VN_out_sig(4919);
CN_in_sig(639)	<=	VN_out_sig(4920);
CN_in_sig(2255)	<=	VN_out_sig(4921);
CN_in_sig(2623)	<=	VN_out_sig(4922);
CN_in_sig(4311)	<=	VN_out_sig(4923);
CN_in_sig(647)	<=	VN_out_sig(4924);
CN_in_sig(2263)	<=	VN_out_sig(4925);
CN_in_sig(2631)	<=	VN_out_sig(4926);
CN_in_sig(4319)	<=	VN_out_sig(4927);
CN_in_sig(655)	<=	VN_out_sig(4928);
CN_in_sig(2271)	<=	VN_out_sig(4929);
CN_in_sig(2639)	<=	VN_out_sig(4930);
CN_in_sig(3895)	<=	VN_out_sig(4931);
CN_in_sig(663)	<=	VN_out_sig(4932);
CN_in_sig(2279)	<=	VN_out_sig(4933);
CN_in_sig(2647)	<=	VN_out_sig(4934);
CN_in_sig(3903)	<=	VN_out_sig(4935);
CN_in_sig(671)	<=	VN_out_sig(4936);
CN_in_sig(2287)	<=	VN_out_sig(4937);
CN_in_sig(2655)	<=	VN_out_sig(4938);
CN_in_sig(3911)	<=	VN_out_sig(4939);
CN_in_sig(679)	<=	VN_out_sig(4940);
CN_in_sig(2295)	<=	VN_out_sig(4941);
CN_in_sig(2663)	<=	VN_out_sig(4942);
CN_in_sig(3919)	<=	VN_out_sig(4943);
CN_in_sig(687)	<=	VN_out_sig(4944);
CN_in_sig(2303)	<=	VN_out_sig(4945);
CN_in_sig(2671)	<=	VN_out_sig(4946);
CN_in_sig(3927)	<=	VN_out_sig(4947);
CN_in_sig(695)	<=	VN_out_sig(4948);
CN_in_sig(2311)	<=	VN_out_sig(4949);
CN_in_sig(2679)	<=	VN_out_sig(4950);
CN_in_sig(3935)	<=	VN_out_sig(4951);
CN_in_sig(703)	<=	VN_out_sig(4952);
CN_in_sig(2319)	<=	VN_out_sig(4953);
CN_in_sig(2687)	<=	VN_out_sig(4954);
CN_in_sig(3943)	<=	VN_out_sig(4955);
CN_in_sig(711)	<=	VN_out_sig(4956);
CN_in_sig(2327)	<=	VN_out_sig(4957);
CN_in_sig(2695)	<=	VN_out_sig(4958);
CN_in_sig(3951)	<=	VN_out_sig(4959);
CN_in_sig(719)	<=	VN_out_sig(4960);
CN_in_sig(2335)	<=	VN_out_sig(4961);
CN_in_sig(2703)	<=	VN_out_sig(4962);
CN_in_sig(3959)	<=	VN_out_sig(4963);
CN_in_sig(727)	<=	VN_out_sig(4964);
CN_in_sig(2343)	<=	VN_out_sig(4965);
CN_in_sig(2711)	<=	VN_out_sig(4966);
CN_in_sig(3967)	<=	VN_out_sig(4967);
CN_in_sig(7)	<=	VN_out_sig(4968);
CN_in_sig(1519)	<=	VN_out_sig(4969);
CN_in_sig(3567)	<=	VN_out_sig(4970);
CN_in_sig(5071)	<=	VN_out_sig(4971);
CN_in_sig(15)	<=	VN_out_sig(4972);
CN_in_sig(1527)	<=	VN_out_sig(4973);
CN_in_sig(3575)	<=	VN_out_sig(4974);
CN_in_sig(5079)	<=	VN_out_sig(4975);
CN_in_sig(23)	<=	VN_out_sig(4976);
CN_in_sig(1535)	<=	VN_out_sig(4977);
CN_in_sig(3583)	<=	VN_out_sig(4978);
CN_in_sig(5087)	<=	VN_out_sig(4979);
CN_in_sig(31)	<=	VN_out_sig(4980);
CN_in_sig(1543)	<=	VN_out_sig(4981);
CN_in_sig(3591)	<=	VN_out_sig(4982);
CN_in_sig(5095)	<=	VN_out_sig(4983);
CN_in_sig(39)	<=	VN_out_sig(4984);
CN_in_sig(1551)	<=	VN_out_sig(4985);
CN_in_sig(3599)	<=	VN_out_sig(4986);
CN_in_sig(5103)	<=	VN_out_sig(4987);
CN_in_sig(47)	<=	VN_out_sig(4988);
CN_in_sig(1559)	<=	VN_out_sig(4989);
CN_in_sig(3607)	<=	VN_out_sig(4990);
CN_in_sig(5111)	<=	VN_out_sig(4991);
CN_in_sig(55)	<=	VN_out_sig(4992);
CN_in_sig(1567)	<=	VN_out_sig(4993);
CN_in_sig(3615)	<=	VN_out_sig(4994);
CN_in_sig(5119)	<=	VN_out_sig(4995);
CN_in_sig(63)	<=	VN_out_sig(4996);
CN_in_sig(1575)	<=	VN_out_sig(4997);
CN_in_sig(3623)	<=	VN_out_sig(4998);
CN_in_sig(5127)	<=	VN_out_sig(4999);
CN_in_sig(71)	<=	VN_out_sig(5000);
CN_in_sig(1583)	<=	VN_out_sig(5001);
CN_in_sig(3631)	<=	VN_out_sig(5002);
CN_in_sig(5135)	<=	VN_out_sig(5003);
CN_in_sig(79)	<=	VN_out_sig(5004);
CN_in_sig(1591)	<=	VN_out_sig(5005);
CN_in_sig(3639)	<=	VN_out_sig(5006);
CN_in_sig(5143)	<=	VN_out_sig(5007);
CN_in_sig(87)	<=	VN_out_sig(5008);
CN_in_sig(1599)	<=	VN_out_sig(5009);
CN_in_sig(3647)	<=	VN_out_sig(5010);
CN_in_sig(5151)	<=	VN_out_sig(5011);
CN_in_sig(95)	<=	VN_out_sig(5012);
CN_in_sig(1607)	<=	VN_out_sig(5013);
CN_in_sig(3655)	<=	VN_out_sig(5014);
CN_in_sig(5159)	<=	VN_out_sig(5015);
CN_in_sig(103)	<=	VN_out_sig(5016);
CN_in_sig(1615)	<=	VN_out_sig(5017);
CN_in_sig(3663)	<=	VN_out_sig(5018);
CN_in_sig(5167)	<=	VN_out_sig(5019);
CN_in_sig(111)	<=	VN_out_sig(5020);
CN_in_sig(1623)	<=	VN_out_sig(5021);
CN_in_sig(3671)	<=	VN_out_sig(5022);
CN_in_sig(5175)	<=	VN_out_sig(5023);
CN_in_sig(119)	<=	VN_out_sig(5024);
CN_in_sig(1631)	<=	VN_out_sig(5025);
CN_in_sig(3679)	<=	VN_out_sig(5026);
CN_in_sig(5183)	<=	VN_out_sig(5027);
CN_in_sig(127)	<=	VN_out_sig(5028);
CN_in_sig(1639)	<=	VN_out_sig(5029);
CN_in_sig(3687)	<=	VN_out_sig(5030);
CN_in_sig(4759)	<=	VN_out_sig(5031);
CN_in_sig(135)	<=	VN_out_sig(5032);
CN_in_sig(1647)	<=	VN_out_sig(5033);
CN_in_sig(3695)	<=	VN_out_sig(5034);
CN_in_sig(4767)	<=	VN_out_sig(5035);
CN_in_sig(143)	<=	VN_out_sig(5036);
CN_in_sig(1655)	<=	VN_out_sig(5037);
CN_in_sig(3703)	<=	VN_out_sig(5038);
CN_in_sig(4775)	<=	VN_out_sig(5039);
CN_in_sig(151)	<=	VN_out_sig(5040);
CN_in_sig(1663)	<=	VN_out_sig(5041);
CN_in_sig(3711)	<=	VN_out_sig(5042);
CN_in_sig(4783)	<=	VN_out_sig(5043);
CN_in_sig(159)	<=	VN_out_sig(5044);
CN_in_sig(1671)	<=	VN_out_sig(5045);
CN_in_sig(3719)	<=	VN_out_sig(5046);
CN_in_sig(4791)	<=	VN_out_sig(5047);
CN_in_sig(167)	<=	VN_out_sig(5048);
CN_in_sig(1679)	<=	VN_out_sig(5049);
CN_in_sig(3727)	<=	VN_out_sig(5050);
CN_in_sig(4799)	<=	VN_out_sig(5051);
CN_in_sig(175)	<=	VN_out_sig(5052);
CN_in_sig(1687)	<=	VN_out_sig(5053);
CN_in_sig(3735)	<=	VN_out_sig(5054);
CN_in_sig(4807)	<=	VN_out_sig(5055);
CN_in_sig(183)	<=	VN_out_sig(5056);
CN_in_sig(1695)	<=	VN_out_sig(5057);
CN_in_sig(3743)	<=	VN_out_sig(5058);
CN_in_sig(4815)	<=	VN_out_sig(5059);
CN_in_sig(191)	<=	VN_out_sig(5060);
CN_in_sig(1703)	<=	VN_out_sig(5061);
CN_in_sig(3751)	<=	VN_out_sig(5062);
CN_in_sig(4823)	<=	VN_out_sig(5063);
CN_in_sig(199)	<=	VN_out_sig(5064);
CN_in_sig(1711)	<=	VN_out_sig(5065);
CN_in_sig(3759)	<=	VN_out_sig(5066);
CN_in_sig(4831)	<=	VN_out_sig(5067);
CN_in_sig(207)	<=	VN_out_sig(5068);
CN_in_sig(1719)	<=	VN_out_sig(5069);
CN_in_sig(3767)	<=	VN_out_sig(5070);
CN_in_sig(4839)	<=	VN_out_sig(5071);
CN_in_sig(215)	<=	VN_out_sig(5072);
CN_in_sig(1727)	<=	VN_out_sig(5073);
CN_in_sig(3775)	<=	VN_out_sig(5074);
CN_in_sig(4847)	<=	VN_out_sig(5075);
CN_in_sig(223)	<=	VN_out_sig(5076);
CN_in_sig(1303)	<=	VN_out_sig(5077);
CN_in_sig(3783)	<=	VN_out_sig(5078);
CN_in_sig(4855)	<=	VN_out_sig(5079);
CN_in_sig(231)	<=	VN_out_sig(5080);
CN_in_sig(1311)	<=	VN_out_sig(5081);
CN_in_sig(3791)	<=	VN_out_sig(5082);
CN_in_sig(4863)	<=	VN_out_sig(5083);
CN_in_sig(239)	<=	VN_out_sig(5084);
CN_in_sig(1319)	<=	VN_out_sig(5085);
CN_in_sig(3799)	<=	VN_out_sig(5086);
CN_in_sig(4871)	<=	VN_out_sig(5087);
CN_in_sig(247)	<=	VN_out_sig(5088);
CN_in_sig(1327)	<=	VN_out_sig(5089);
CN_in_sig(3807)	<=	VN_out_sig(5090);
CN_in_sig(4879)	<=	VN_out_sig(5091);
CN_in_sig(255)	<=	VN_out_sig(5092);
CN_in_sig(1335)	<=	VN_out_sig(5093);
CN_in_sig(3815)	<=	VN_out_sig(5094);
CN_in_sig(4887)	<=	VN_out_sig(5095);
CN_in_sig(263)	<=	VN_out_sig(5096);
CN_in_sig(1343)	<=	VN_out_sig(5097);
CN_in_sig(3823)	<=	VN_out_sig(5098);
CN_in_sig(4895)	<=	VN_out_sig(5099);
CN_in_sig(271)	<=	VN_out_sig(5100);
CN_in_sig(1351)	<=	VN_out_sig(5101);
CN_in_sig(3831)	<=	VN_out_sig(5102);
CN_in_sig(4903)	<=	VN_out_sig(5103);
CN_in_sig(279)	<=	VN_out_sig(5104);
CN_in_sig(1359)	<=	VN_out_sig(5105);
CN_in_sig(3839)	<=	VN_out_sig(5106);
CN_in_sig(4911)	<=	VN_out_sig(5107);
CN_in_sig(287)	<=	VN_out_sig(5108);
CN_in_sig(1367)	<=	VN_out_sig(5109);
CN_in_sig(3847)	<=	VN_out_sig(5110);
CN_in_sig(4919)	<=	VN_out_sig(5111);
CN_in_sig(295)	<=	VN_out_sig(5112);
CN_in_sig(1375)	<=	VN_out_sig(5113);
CN_in_sig(3855)	<=	VN_out_sig(5114);
CN_in_sig(4927)	<=	VN_out_sig(5115);
CN_in_sig(303)	<=	VN_out_sig(5116);
CN_in_sig(1383)	<=	VN_out_sig(5117);
CN_in_sig(3863)	<=	VN_out_sig(5118);
CN_in_sig(4935)	<=	VN_out_sig(5119);
CN_in_sig(311)	<=	VN_out_sig(5120);
CN_in_sig(1391)	<=	VN_out_sig(5121);
CN_in_sig(3871)	<=	VN_out_sig(5122);
CN_in_sig(4943)	<=	VN_out_sig(5123);
CN_in_sig(319)	<=	VN_out_sig(5124);
CN_in_sig(1399)	<=	VN_out_sig(5125);
CN_in_sig(3879)	<=	VN_out_sig(5126);
CN_in_sig(4951)	<=	VN_out_sig(5127);
CN_in_sig(327)	<=	VN_out_sig(5128);
CN_in_sig(1407)	<=	VN_out_sig(5129);
CN_in_sig(3887)	<=	VN_out_sig(5130);
CN_in_sig(4959)	<=	VN_out_sig(5131);
CN_in_sig(335)	<=	VN_out_sig(5132);
CN_in_sig(1415)	<=	VN_out_sig(5133);
CN_in_sig(3463)	<=	VN_out_sig(5134);
CN_in_sig(4967)	<=	VN_out_sig(5135);
CN_in_sig(343)	<=	VN_out_sig(5136);
CN_in_sig(1423)	<=	VN_out_sig(5137);
CN_in_sig(3471)	<=	VN_out_sig(5138);
CN_in_sig(4975)	<=	VN_out_sig(5139);
CN_in_sig(351)	<=	VN_out_sig(5140);
CN_in_sig(1431)	<=	VN_out_sig(5141);
CN_in_sig(3479)	<=	VN_out_sig(5142);
CN_in_sig(4983)	<=	VN_out_sig(5143);
CN_in_sig(359)	<=	VN_out_sig(5144);
CN_in_sig(1439)	<=	VN_out_sig(5145);
CN_in_sig(3487)	<=	VN_out_sig(5146);
CN_in_sig(4991)	<=	VN_out_sig(5147);
CN_in_sig(367)	<=	VN_out_sig(5148);
CN_in_sig(1447)	<=	VN_out_sig(5149);
CN_in_sig(3495)	<=	VN_out_sig(5150);
CN_in_sig(4999)	<=	VN_out_sig(5151);
CN_in_sig(375)	<=	VN_out_sig(5152);
CN_in_sig(1455)	<=	VN_out_sig(5153);
CN_in_sig(3503)	<=	VN_out_sig(5154);
CN_in_sig(5007)	<=	VN_out_sig(5155);
CN_in_sig(383)	<=	VN_out_sig(5156);
CN_in_sig(1463)	<=	VN_out_sig(5157);
CN_in_sig(3511)	<=	VN_out_sig(5158);
CN_in_sig(5015)	<=	VN_out_sig(5159);
CN_in_sig(391)	<=	VN_out_sig(5160);
CN_in_sig(1471)	<=	VN_out_sig(5161);
CN_in_sig(3519)	<=	VN_out_sig(5162);
CN_in_sig(5023)	<=	VN_out_sig(5163);
CN_in_sig(399)	<=	VN_out_sig(5164);
CN_in_sig(1479)	<=	VN_out_sig(5165);
CN_in_sig(3527)	<=	VN_out_sig(5166);
CN_in_sig(5031)	<=	VN_out_sig(5167);
CN_in_sig(407)	<=	VN_out_sig(5168);
CN_in_sig(1487)	<=	VN_out_sig(5169);
CN_in_sig(3535)	<=	VN_out_sig(5170);
CN_in_sig(5039)	<=	VN_out_sig(5171);
CN_in_sig(415)	<=	VN_out_sig(5172);
CN_in_sig(1495)	<=	VN_out_sig(5173);
CN_in_sig(3543)	<=	VN_out_sig(5174);
CN_in_sig(5047)	<=	VN_out_sig(5175);
CN_in_sig(423)	<=	VN_out_sig(5176);
CN_in_sig(1503)	<=	VN_out_sig(5177);
CN_in_sig(3551)	<=	VN_out_sig(5178);
CN_in_sig(5055)	<=	VN_out_sig(5179);
CN_in_sig(431)	<=	VN_out_sig(5180);
CN_in_sig(1511)	<=	VN_out_sig(5181);
CN_in_sig(3559)	<=	VN_out_sig(5182);
CN_in_sig(5063)	<=	VN_out_sig(5183);


CN_in_sigd(344)	<=	VN_out_sigd(0);
CN_in_sigd(1512)	<=	VN_out_sigd(0);
CN_in_sigd(3816)	<=	VN_out_sigd(0);
CN_in_sigd(4872)	<=	VN_out_sigd(0);
CN_in_sigd(352)	<=	VN_out_sigd(1);
CN_in_sigd(1520)	<=	VN_out_sigd(1);
CN_in_sigd(3824)	<=	VN_out_sigd(1);
CN_in_sigd(4880)	<=	VN_out_sigd(1);
CN_in_sigd(360)	<=	VN_out_sigd(2);
CN_in_sigd(1528)	<=	VN_out_sigd(2);
CN_in_sigd(3832)	<=	VN_out_sigd(2);
CN_in_sigd(4888)	<=	VN_out_sigd(2);
CN_in_sigd(368)	<=	VN_out_sigd(3);
CN_in_sigd(1536)	<=	VN_out_sigd(3);
CN_in_sigd(3840)	<=	VN_out_sigd(3);
CN_in_sigd(4896)	<=	VN_out_sigd(3);
CN_in_sigd(376)	<=	VN_out_sigd(4);
CN_in_sigd(1544)	<=	VN_out_sigd(4);
CN_in_sigd(3848)	<=	VN_out_sigd(4);
CN_in_sigd(4904)	<=	VN_out_sigd(4);
CN_in_sigd(384)	<=	VN_out_sigd(5);
CN_in_sigd(1552)	<=	VN_out_sigd(5);
CN_in_sigd(3856)	<=	VN_out_sigd(5);
CN_in_sigd(4912)	<=	VN_out_sigd(5);
CN_in_sigd(392)	<=	VN_out_sigd(6);
CN_in_sigd(1560)	<=	VN_out_sigd(6);
CN_in_sigd(3864)	<=	VN_out_sigd(6);
CN_in_sigd(4920)	<=	VN_out_sigd(6);
CN_in_sigd(400)	<=	VN_out_sigd(7);
CN_in_sigd(1568)	<=	VN_out_sigd(7);
CN_in_sigd(3872)	<=	VN_out_sigd(7);
CN_in_sigd(4928)	<=	VN_out_sigd(7);
CN_in_sigd(408)	<=	VN_out_sigd(8);
CN_in_sigd(1576)	<=	VN_out_sigd(8);
CN_in_sigd(3880)	<=	VN_out_sigd(8);
CN_in_sigd(4936)	<=	VN_out_sigd(8);
CN_in_sigd(416)	<=	VN_out_sigd(9);
CN_in_sigd(1584)	<=	VN_out_sigd(9);
CN_in_sigd(3456)	<=	VN_out_sigd(9);
CN_in_sigd(4944)	<=	VN_out_sigd(9);
CN_in_sigd(424)	<=	VN_out_sigd(10);
CN_in_sigd(1592)	<=	VN_out_sigd(10);
CN_in_sigd(3464)	<=	VN_out_sigd(10);
CN_in_sigd(4952)	<=	VN_out_sigd(10);
CN_in_sigd(0)	<=	VN_out_sigd(11);
CN_in_sigd(1600)	<=	VN_out_sigd(11);
CN_in_sigd(3472)	<=	VN_out_sigd(11);
CN_in_sigd(4960)	<=	VN_out_sigd(11);
CN_in_sigd(8)	<=	VN_out_sigd(12);
CN_in_sigd(1608)	<=	VN_out_sigd(12);
CN_in_sigd(3480)	<=	VN_out_sigd(12);
CN_in_sigd(4968)	<=	VN_out_sigd(12);
CN_in_sigd(16)	<=	VN_out_sigd(13);
CN_in_sigd(1616)	<=	VN_out_sigd(13);
CN_in_sigd(3488)	<=	VN_out_sigd(13);
CN_in_sigd(4976)	<=	VN_out_sigd(13);
CN_in_sigd(24)	<=	VN_out_sigd(14);
CN_in_sigd(1624)	<=	VN_out_sigd(14);
CN_in_sigd(3496)	<=	VN_out_sigd(14);
CN_in_sigd(4984)	<=	VN_out_sigd(14);
CN_in_sigd(32)	<=	VN_out_sigd(15);
CN_in_sigd(1632)	<=	VN_out_sigd(15);
CN_in_sigd(3504)	<=	VN_out_sigd(15);
CN_in_sigd(4992)	<=	VN_out_sigd(15);
CN_in_sigd(40)	<=	VN_out_sigd(16);
CN_in_sigd(1640)	<=	VN_out_sigd(16);
CN_in_sigd(3512)	<=	VN_out_sigd(16);
CN_in_sigd(5000)	<=	VN_out_sigd(16);
CN_in_sigd(48)	<=	VN_out_sigd(17);
CN_in_sigd(1648)	<=	VN_out_sigd(17);
CN_in_sigd(3520)	<=	VN_out_sigd(17);
CN_in_sigd(5008)	<=	VN_out_sigd(17);
CN_in_sigd(56)	<=	VN_out_sigd(18);
CN_in_sigd(1656)	<=	VN_out_sigd(18);
CN_in_sigd(3528)	<=	VN_out_sigd(18);
CN_in_sigd(5016)	<=	VN_out_sigd(18);
CN_in_sigd(64)	<=	VN_out_sigd(19);
CN_in_sigd(1664)	<=	VN_out_sigd(19);
CN_in_sigd(3536)	<=	VN_out_sigd(19);
CN_in_sigd(5024)	<=	VN_out_sigd(19);
CN_in_sigd(72)	<=	VN_out_sigd(20);
CN_in_sigd(1672)	<=	VN_out_sigd(20);
CN_in_sigd(3544)	<=	VN_out_sigd(20);
CN_in_sigd(5032)	<=	VN_out_sigd(20);
CN_in_sigd(80)	<=	VN_out_sigd(21);
CN_in_sigd(1680)	<=	VN_out_sigd(21);
CN_in_sigd(3552)	<=	VN_out_sigd(21);
CN_in_sigd(5040)	<=	VN_out_sigd(21);
CN_in_sigd(88)	<=	VN_out_sigd(22);
CN_in_sigd(1688)	<=	VN_out_sigd(22);
CN_in_sigd(3560)	<=	VN_out_sigd(22);
CN_in_sigd(5048)	<=	VN_out_sigd(22);
CN_in_sigd(96)	<=	VN_out_sigd(23);
CN_in_sigd(1696)	<=	VN_out_sigd(23);
CN_in_sigd(3568)	<=	VN_out_sigd(23);
CN_in_sigd(5056)	<=	VN_out_sigd(23);
CN_in_sigd(104)	<=	VN_out_sigd(24);
CN_in_sigd(1704)	<=	VN_out_sigd(24);
CN_in_sigd(3576)	<=	VN_out_sigd(24);
CN_in_sigd(5064)	<=	VN_out_sigd(24);
CN_in_sigd(112)	<=	VN_out_sigd(25);
CN_in_sigd(1712)	<=	VN_out_sigd(25);
CN_in_sigd(3584)	<=	VN_out_sigd(25);
CN_in_sigd(5072)	<=	VN_out_sigd(25);
CN_in_sigd(120)	<=	VN_out_sigd(26);
CN_in_sigd(1720)	<=	VN_out_sigd(26);
CN_in_sigd(3592)	<=	VN_out_sigd(26);
CN_in_sigd(5080)	<=	VN_out_sigd(26);
CN_in_sigd(128)	<=	VN_out_sigd(27);
CN_in_sigd(1296)	<=	VN_out_sigd(27);
CN_in_sigd(3600)	<=	VN_out_sigd(27);
CN_in_sigd(5088)	<=	VN_out_sigd(27);
CN_in_sigd(136)	<=	VN_out_sigd(28);
CN_in_sigd(1304)	<=	VN_out_sigd(28);
CN_in_sigd(3608)	<=	VN_out_sigd(28);
CN_in_sigd(5096)	<=	VN_out_sigd(28);
CN_in_sigd(144)	<=	VN_out_sigd(29);
CN_in_sigd(1312)	<=	VN_out_sigd(29);
CN_in_sigd(3616)	<=	VN_out_sigd(29);
CN_in_sigd(5104)	<=	VN_out_sigd(29);
CN_in_sigd(152)	<=	VN_out_sigd(30);
CN_in_sigd(1320)	<=	VN_out_sigd(30);
CN_in_sigd(3624)	<=	VN_out_sigd(30);
CN_in_sigd(5112)	<=	VN_out_sigd(30);
CN_in_sigd(160)	<=	VN_out_sigd(31);
CN_in_sigd(1328)	<=	VN_out_sigd(31);
CN_in_sigd(3632)	<=	VN_out_sigd(31);
CN_in_sigd(5120)	<=	VN_out_sigd(31);
CN_in_sigd(168)	<=	VN_out_sigd(32);
CN_in_sigd(1336)	<=	VN_out_sigd(32);
CN_in_sigd(3640)	<=	VN_out_sigd(32);
CN_in_sigd(5128)	<=	VN_out_sigd(32);
CN_in_sigd(176)	<=	VN_out_sigd(33);
CN_in_sigd(1344)	<=	VN_out_sigd(33);
CN_in_sigd(3648)	<=	VN_out_sigd(33);
CN_in_sigd(5136)	<=	VN_out_sigd(33);
CN_in_sigd(184)	<=	VN_out_sigd(34);
CN_in_sigd(1352)	<=	VN_out_sigd(34);
CN_in_sigd(3656)	<=	VN_out_sigd(34);
CN_in_sigd(5144)	<=	VN_out_sigd(34);
CN_in_sigd(192)	<=	VN_out_sigd(35);
CN_in_sigd(1360)	<=	VN_out_sigd(35);
CN_in_sigd(3664)	<=	VN_out_sigd(35);
CN_in_sigd(5152)	<=	VN_out_sigd(35);
CN_in_sigd(200)	<=	VN_out_sigd(36);
CN_in_sigd(1368)	<=	VN_out_sigd(36);
CN_in_sigd(3672)	<=	VN_out_sigd(36);
CN_in_sigd(5160)	<=	VN_out_sigd(36);
CN_in_sigd(208)	<=	VN_out_sigd(37);
CN_in_sigd(1376)	<=	VN_out_sigd(37);
CN_in_sigd(3680)	<=	VN_out_sigd(37);
CN_in_sigd(5168)	<=	VN_out_sigd(37);
CN_in_sigd(216)	<=	VN_out_sigd(38);
CN_in_sigd(1384)	<=	VN_out_sigd(38);
CN_in_sigd(3688)	<=	VN_out_sigd(38);
CN_in_sigd(5176)	<=	VN_out_sigd(38);
CN_in_sigd(224)	<=	VN_out_sigd(39);
CN_in_sigd(1392)	<=	VN_out_sigd(39);
CN_in_sigd(3696)	<=	VN_out_sigd(39);
CN_in_sigd(4752)	<=	VN_out_sigd(39);
CN_in_sigd(232)	<=	VN_out_sigd(40);
CN_in_sigd(1400)	<=	VN_out_sigd(40);
CN_in_sigd(3704)	<=	VN_out_sigd(40);
CN_in_sigd(4760)	<=	VN_out_sigd(40);
CN_in_sigd(240)	<=	VN_out_sigd(41);
CN_in_sigd(1408)	<=	VN_out_sigd(41);
CN_in_sigd(3712)	<=	VN_out_sigd(41);
CN_in_sigd(4768)	<=	VN_out_sigd(41);
CN_in_sigd(248)	<=	VN_out_sigd(42);
CN_in_sigd(1416)	<=	VN_out_sigd(42);
CN_in_sigd(3720)	<=	VN_out_sigd(42);
CN_in_sigd(4776)	<=	VN_out_sigd(42);
CN_in_sigd(256)	<=	VN_out_sigd(43);
CN_in_sigd(1424)	<=	VN_out_sigd(43);
CN_in_sigd(3728)	<=	VN_out_sigd(43);
CN_in_sigd(4784)	<=	VN_out_sigd(43);
CN_in_sigd(264)	<=	VN_out_sigd(44);
CN_in_sigd(1432)	<=	VN_out_sigd(44);
CN_in_sigd(3736)	<=	VN_out_sigd(44);
CN_in_sigd(4792)	<=	VN_out_sigd(44);
CN_in_sigd(272)	<=	VN_out_sigd(45);
CN_in_sigd(1440)	<=	VN_out_sigd(45);
CN_in_sigd(3744)	<=	VN_out_sigd(45);
CN_in_sigd(4800)	<=	VN_out_sigd(45);
CN_in_sigd(280)	<=	VN_out_sigd(46);
CN_in_sigd(1448)	<=	VN_out_sigd(46);
CN_in_sigd(3752)	<=	VN_out_sigd(46);
CN_in_sigd(4808)	<=	VN_out_sigd(46);
CN_in_sigd(288)	<=	VN_out_sigd(47);
CN_in_sigd(1456)	<=	VN_out_sigd(47);
CN_in_sigd(3760)	<=	VN_out_sigd(47);
CN_in_sigd(4816)	<=	VN_out_sigd(47);
CN_in_sigd(296)	<=	VN_out_sigd(48);
CN_in_sigd(1464)	<=	VN_out_sigd(48);
CN_in_sigd(3768)	<=	VN_out_sigd(48);
CN_in_sigd(4824)	<=	VN_out_sigd(48);
CN_in_sigd(304)	<=	VN_out_sigd(49);
CN_in_sigd(1472)	<=	VN_out_sigd(49);
CN_in_sigd(3776)	<=	VN_out_sigd(49);
CN_in_sigd(4832)	<=	VN_out_sigd(49);
CN_in_sigd(312)	<=	VN_out_sigd(50);
CN_in_sigd(1480)	<=	VN_out_sigd(50);
CN_in_sigd(3784)	<=	VN_out_sigd(50);
CN_in_sigd(4840)	<=	VN_out_sigd(50);
CN_in_sigd(320)	<=	VN_out_sigd(51);
CN_in_sigd(1488)	<=	VN_out_sigd(51);
CN_in_sigd(3792)	<=	VN_out_sigd(51);
CN_in_sigd(4848)	<=	VN_out_sigd(51);
CN_in_sigd(328)	<=	VN_out_sigd(52);
CN_in_sigd(1496)	<=	VN_out_sigd(52);
CN_in_sigd(3800)	<=	VN_out_sigd(52);
CN_in_sigd(4856)	<=	VN_out_sigd(52);
CN_in_sigd(336)	<=	VN_out_sigd(53);
CN_in_sigd(1504)	<=	VN_out_sigd(53);
CN_in_sigd(3808)	<=	VN_out_sigd(53);
CN_in_sigd(4864)	<=	VN_out_sigd(53);
CN_in_sigd(664)	<=	VN_out_sigd(54);
CN_in_sigd(1824)	<=	VN_out_sigd(54);
CN_in_sigd(3224)	<=	VN_out_sigd(54);
CN_in_sigd(4720)	<=	VN_out_sigd(54);
CN_in_sigd(672)	<=	VN_out_sigd(55);
CN_in_sigd(1832)	<=	VN_out_sigd(55);
CN_in_sigd(3232)	<=	VN_out_sigd(55);
CN_in_sigd(4728)	<=	VN_out_sigd(55);
CN_in_sigd(680)	<=	VN_out_sigd(56);
CN_in_sigd(1840)	<=	VN_out_sigd(56);
CN_in_sigd(3240)	<=	VN_out_sigd(56);
CN_in_sigd(4736)	<=	VN_out_sigd(56);
CN_in_sigd(688)	<=	VN_out_sigd(57);
CN_in_sigd(1848)	<=	VN_out_sigd(57);
CN_in_sigd(3248)	<=	VN_out_sigd(57);
CN_in_sigd(4744)	<=	VN_out_sigd(57);
CN_in_sigd(696)	<=	VN_out_sigd(58);
CN_in_sigd(1856)	<=	VN_out_sigd(58);
CN_in_sigd(3256)	<=	VN_out_sigd(58);
CN_in_sigd(4320)	<=	VN_out_sigd(58);
CN_in_sigd(704)	<=	VN_out_sigd(59);
CN_in_sigd(1864)	<=	VN_out_sigd(59);
CN_in_sigd(3264)	<=	VN_out_sigd(59);
CN_in_sigd(4328)	<=	VN_out_sigd(59);
CN_in_sigd(712)	<=	VN_out_sigd(60);
CN_in_sigd(1872)	<=	VN_out_sigd(60);
CN_in_sigd(3272)	<=	VN_out_sigd(60);
CN_in_sigd(4336)	<=	VN_out_sigd(60);
CN_in_sigd(720)	<=	VN_out_sigd(61);
CN_in_sigd(1880)	<=	VN_out_sigd(61);
CN_in_sigd(3280)	<=	VN_out_sigd(61);
CN_in_sigd(4344)	<=	VN_out_sigd(61);
CN_in_sigd(728)	<=	VN_out_sigd(62);
CN_in_sigd(1888)	<=	VN_out_sigd(62);
CN_in_sigd(3288)	<=	VN_out_sigd(62);
CN_in_sigd(4352)	<=	VN_out_sigd(62);
CN_in_sigd(736)	<=	VN_out_sigd(63);
CN_in_sigd(1896)	<=	VN_out_sigd(63);
CN_in_sigd(3296)	<=	VN_out_sigd(63);
CN_in_sigd(4360)	<=	VN_out_sigd(63);
CN_in_sigd(744)	<=	VN_out_sigd(64);
CN_in_sigd(1904)	<=	VN_out_sigd(64);
CN_in_sigd(3304)	<=	VN_out_sigd(64);
CN_in_sigd(4368)	<=	VN_out_sigd(64);
CN_in_sigd(752)	<=	VN_out_sigd(65);
CN_in_sigd(1912)	<=	VN_out_sigd(65);
CN_in_sigd(3312)	<=	VN_out_sigd(65);
CN_in_sigd(4376)	<=	VN_out_sigd(65);
CN_in_sigd(760)	<=	VN_out_sigd(66);
CN_in_sigd(1920)	<=	VN_out_sigd(66);
CN_in_sigd(3320)	<=	VN_out_sigd(66);
CN_in_sigd(4384)	<=	VN_out_sigd(66);
CN_in_sigd(768)	<=	VN_out_sigd(67);
CN_in_sigd(1928)	<=	VN_out_sigd(67);
CN_in_sigd(3328)	<=	VN_out_sigd(67);
CN_in_sigd(4392)	<=	VN_out_sigd(67);
CN_in_sigd(776)	<=	VN_out_sigd(68);
CN_in_sigd(1936)	<=	VN_out_sigd(68);
CN_in_sigd(3336)	<=	VN_out_sigd(68);
CN_in_sigd(4400)	<=	VN_out_sigd(68);
CN_in_sigd(784)	<=	VN_out_sigd(69);
CN_in_sigd(1944)	<=	VN_out_sigd(69);
CN_in_sigd(3344)	<=	VN_out_sigd(69);
CN_in_sigd(4408)	<=	VN_out_sigd(69);
CN_in_sigd(792)	<=	VN_out_sigd(70);
CN_in_sigd(1952)	<=	VN_out_sigd(70);
CN_in_sigd(3352)	<=	VN_out_sigd(70);
CN_in_sigd(4416)	<=	VN_out_sigd(70);
CN_in_sigd(800)	<=	VN_out_sigd(71);
CN_in_sigd(1960)	<=	VN_out_sigd(71);
CN_in_sigd(3360)	<=	VN_out_sigd(71);
CN_in_sigd(4424)	<=	VN_out_sigd(71);
CN_in_sigd(808)	<=	VN_out_sigd(72);
CN_in_sigd(1968)	<=	VN_out_sigd(72);
CN_in_sigd(3368)	<=	VN_out_sigd(72);
CN_in_sigd(4432)	<=	VN_out_sigd(72);
CN_in_sigd(816)	<=	VN_out_sigd(73);
CN_in_sigd(1976)	<=	VN_out_sigd(73);
CN_in_sigd(3376)	<=	VN_out_sigd(73);
CN_in_sigd(4440)	<=	VN_out_sigd(73);
CN_in_sigd(824)	<=	VN_out_sigd(74);
CN_in_sigd(1984)	<=	VN_out_sigd(74);
CN_in_sigd(3384)	<=	VN_out_sigd(74);
CN_in_sigd(4448)	<=	VN_out_sigd(74);
CN_in_sigd(832)	<=	VN_out_sigd(75);
CN_in_sigd(1992)	<=	VN_out_sigd(75);
CN_in_sigd(3392)	<=	VN_out_sigd(75);
CN_in_sigd(4456)	<=	VN_out_sigd(75);
CN_in_sigd(840)	<=	VN_out_sigd(76);
CN_in_sigd(2000)	<=	VN_out_sigd(76);
CN_in_sigd(3400)	<=	VN_out_sigd(76);
CN_in_sigd(4464)	<=	VN_out_sigd(76);
CN_in_sigd(848)	<=	VN_out_sigd(77);
CN_in_sigd(2008)	<=	VN_out_sigd(77);
CN_in_sigd(3408)	<=	VN_out_sigd(77);
CN_in_sigd(4472)	<=	VN_out_sigd(77);
CN_in_sigd(856)	<=	VN_out_sigd(78);
CN_in_sigd(2016)	<=	VN_out_sigd(78);
CN_in_sigd(3416)	<=	VN_out_sigd(78);
CN_in_sigd(4480)	<=	VN_out_sigd(78);
CN_in_sigd(432)	<=	VN_out_sigd(79);
CN_in_sigd(2024)	<=	VN_out_sigd(79);
CN_in_sigd(3424)	<=	VN_out_sigd(79);
CN_in_sigd(4488)	<=	VN_out_sigd(79);
CN_in_sigd(440)	<=	VN_out_sigd(80);
CN_in_sigd(2032)	<=	VN_out_sigd(80);
CN_in_sigd(3432)	<=	VN_out_sigd(80);
CN_in_sigd(4496)	<=	VN_out_sigd(80);
CN_in_sigd(448)	<=	VN_out_sigd(81);
CN_in_sigd(2040)	<=	VN_out_sigd(81);
CN_in_sigd(3440)	<=	VN_out_sigd(81);
CN_in_sigd(4504)	<=	VN_out_sigd(81);
CN_in_sigd(456)	<=	VN_out_sigd(82);
CN_in_sigd(2048)	<=	VN_out_sigd(82);
CN_in_sigd(3448)	<=	VN_out_sigd(82);
CN_in_sigd(4512)	<=	VN_out_sigd(82);
CN_in_sigd(464)	<=	VN_out_sigd(83);
CN_in_sigd(2056)	<=	VN_out_sigd(83);
CN_in_sigd(3024)	<=	VN_out_sigd(83);
CN_in_sigd(4520)	<=	VN_out_sigd(83);
CN_in_sigd(472)	<=	VN_out_sigd(84);
CN_in_sigd(2064)	<=	VN_out_sigd(84);
CN_in_sigd(3032)	<=	VN_out_sigd(84);
CN_in_sigd(4528)	<=	VN_out_sigd(84);
CN_in_sigd(480)	<=	VN_out_sigd(85);
CN_in_sigd(2072)	<=	VN_out_sigd(85);
CN_in_sigd(3040)	<=	VN_out_sigd(85);
CN_in_sigd(4536)	<=	VN_out_sigd(85);
CN_in_sigd(488)	<=	VN_out_sigd(86);
CN_in_sigd(2080)	<=	VN_out_sigd(86);
CN_in_sigd(3048)	<=	VN_out_sigd(86);
CN_in_sigd(4544)	<=	VN_out_sigd(86);
CN_in_sigd(496)	<=	VN_out_sigd(87);
CN_in_sigd(2088)	<=	VN_out_sigd(87);
CN_in_sigd(3056)	<=	VN_out_sigd(87);
CN_in_sigd(4552)	<=	VN_out_sigd(87);
CN_in_sigd(504)	<=	VN_out_sigd(88);
CN_in_sigd(2096)	<=	VN_out_sigd(88);
CN_in_sigd(3064)	<=	VN_out_sigd(88);
CN_in_sigd(4560)	<=	VN_out_sigd(88);
CN_in_sigd(512)	<=	VN_out_sigd(89);
CN_in_sigd(2104)	<=	VN_out_sigd(89);
CN_in_sigd(3072)	<=	VN_out_sigd(89);
CN_in_sigd(4568)	<=	VN_out_sigd(89);
CN_in_sigd(520)	<=	VN_out_sigd(90);
CN_in_sigd(2112)	<=	VN_out_sigd(90);
CN_in_sigd(3080)	<=	VN_out_sigd(90);
CN_in_sigd(4576)	<=	VN_out_sigd(90);
CN_in_sigd(528)	<=	VN_out_sigd(91);
CN_in_sigd(2120)	<=	VN_out_sigd(91);
CN_in_sigd(3088)	<=	VN_out_sigd(91);
CN_in_sigd(4584)	<=	VN_out_sigd(91);
CN_in_sigd(536)	<=	VN_out_sigd(92);
CN_in_sigd(2128)	<=	VN_out_sigd(92);
CN_in_sigd(3096)	<=	VN_out_sigd(92);
CN_in_sigd(4592)	<=	VN_out_sigd(92);
CN_in_sigd(544)	<=	VN_out_sigd(93);
CN_in_sigd(2136)	<=	VN_out_sigd(93);
CN_in_sigd(3104)	<=	VN_out_sigd(93);
CN_in_sigd(4600)	<=	VN_out_sigd(93);
CN_in_sigd(552)	<=	VN_out_sigd(94);
CN_in_sigd(2144)	<=	VN_out_sigd(94);
CN_in_sigd(3112)	<=	VN_out_sigd(94);
CN_in_sigd(4608)	<=	VN_out_sigd(94);
CN_in_sigd(560)	<=	VN_out_sigd(95);
CN_in_sigd(2152)	<=	VN_out_sigd(95);
CN_in_sigd(3120)	<=	VN_out_sigd(95);
CN_in_sigd(4616)	<=	VN_out_sigd(95);
CN_in_sigd(568)	<=	VN_out_sigd(96);
CN_in_sigd(1728)	<=	VN_out_sigd(96);
CN_in_sigd(3128)	<=	VN_out_sigd(96);
CN_in_sigd(4624)	<=	VN_out_sigd(96);
CN_in_sigd(576)	<=	VN_out_sigd(97);
CN_in_sigd(1736)	<=	VN_out_sigd(97);
CN_in_sigd(3136)	<=	VN_out_sigd(97);
CN_in_sigd(4632)	<=	VN_out_sigd(97);
CN_in_sigd(584)	<=	VN_out_sigd(98);
CN_in_sigd(1744)	<=	VN_out_sigd(98);
CN_in_sigd(3144)	<=	VN_out_sigd(98);
CN_in_sigd(4640)	<=	VN_out_sigd(98);
CN_in_sigd(592)	<=	VN_out_sigd(99);
CN_in_sigd(1752)	<=	VN_out_sigd(99);
CN_in_sigd(3152)	<=	VN_out_sigd(99);
CN_in_sigd(4648)	<=	VN_out_sigd(99);
CN_in_sigd(600)	<=	VN_out_sigd(100);
CN_in_sigd(1760)	<=	VN_out_sigd(100);
CN_in_sigd(3160)	<=	VN_out_sigd(100);
CN_in_sigd(4656)	<=	VN_out_sigd(100);
CN_in_sigd(608)	<=	VN_out_sigd(101);
CN_in_sigd(1768)	<=	VN_out_sigd(101);
CN_in_sigd(3168)	<=	VN_out_sigd(101);
CN_in_sigd(4664)	<=	VN_out_sigd(101);
CN_in_sigd(616)	<=	VN_out_sigd(102);
CN_in_sigd(1776)	<=	VN_out_sigd(102);
CN_in_sigd(3176)	<=	VN_out_sigd(102);
CN_in_sigd(4672)	<=	VN_out_sigd(102);
CN_in_sigd(624)	<=	VN_out_sigd(103);
CN_in_sigd(1784)	<=	VN_out_sigd(103);
CN_in_sigd(3184)	<=	VN_out_sigd(103);
CN_in_sigd(4680)	<=	VN_out_sigd(103);
CN_in_sigd(632)	<=	VN_out_sigd(104);
CN_in_sigd(1792)	<=	VN_out_sigd(104);
CN_in_sigd(3192)	<=	VN_out_sigd(104);
CN_in_sigd(4688)	<=	VN_out_sigd(104);
CN_in_sigd(640)	<=	VN_out_sigd(105);
CN_in_sigd(1800)	<=	VN_out_sigd(105);
CN_in_sigd(3200)	<=	VN_out_sigd(105);
CN_in_sigd(4696)	<=	VN_out_sigd(105);
CN_in_sigd(648)	<=	VN_out_sigd(106);
CN_in_sigd(1808)	<=	VN_out_sigd(106);
CN_in_sigd(3208)	<=	VN_out_sigd(106);
CN_in_sigd(4704)	<=	VN_out_sigd(106);
CN_in_sigd(656)	<=	VN_out_sigd(107);
CN_in_sigd(1816)	<=	VN_out_sigd(107);
CN_in_sigd(3216)	<=	VN_out_sigd(107);
CN_in_sigd(4712)	<=	VN_out_sigd(107);
CN_in_sigd(944)	<=	VN_out_sigd(108);
CN_in_sigd(2400)	<=	VN_out_sigd(108);
CN_in_sigd(2704)	<=	VN_out_sigd(108);
CN_in_sigd(3896)	<=	VN_out_sigd(108);
CN_in_sigd(952)	<=	VN_out_sigd(109);
CN_in_sigd(2408)	<=	VN_out_sigd(109);
CN_in_sigd(2712)	<=	VN_out_sigd(109);
CN_in_sigd(3904)	<=	VN_out_sigd(109);
CN_in_sigd(960)	<=	VN_out_sigd(110);
CN_in_sigd(2416)	<=	VN_out_sigd(110);
CN_in_sigd(2720)	<=	VN_out_sigd(110);
CN_in_sigd(3912)	<=	VN_out_sigd(110);
CN_in_sigd(968)	<=	VN_out_sigd(111);
CN_in_sigd(2424)	<=	VN_out_sigd(111);
CN_in_sigd(2728)	<=	VN_out_sigd(111);
CN_in_sigd(3920)	<=	VN_out_sigd(111);
CN_in_sigd(976)	<=	VN_out_sigd(112);
CN_in_sigd(2432)	<=	VN_out_sigd(112);
CN_in_sigd(2736)	<=	VN_out_sigd(112);
CN_in_sigd(3928)	<=	VN_out_sigd(112);
CN_in_sigd(984)	<=	VN_out_sigd(113);
CN_in_sigd(2440)	<=	VN_out_sigd(113);
CN_in_sigd(2744)	<=	VN_out_sigd(113);
CN_in_sigd(3936)	<=	VN_out_sigd(113);
CN_in_sigd(992)	<=	VN_out_sigd(114);
CN_in_sigd(2448)	<=	VN_out_sigd(114);
CN_in_sigd(2752)	<=	VN_out_sigd(114);
CN_in_sigd(3944)	<=	VN_out_sigd(114);
CN_in_sigd(1000)	<=	VN_out_sigd(115);
CN_in_sigd(2456)	<=	VN_out_sigd(115);
CN_in_sigd(2760)	<=	VN_out_sigd(115);
CN_in_sigd(3952)	<=	VN_out_sigd(115);
CN_in_sigd(1008)	<=	VN_out_sigd(116);
CN_in_sigd(2464)	<=	VN_out_sigd(116);
CN_in_sigd(2768)	<=	VN_out_sigd(116);
CN_in_sigd(3960)	<=	VN_out_sigd(116);
CN_in_sigd(1016)	<=	VN_out_sigd(117);
CN_in_sigd(2472)	<=	VN_out_sigd(117);
CN_in_sigd(2776)	<=	VN_out_sigd(117);
CN_in_sigd(3968)	<=	VN_out_sigd(117);
CN_in_sigd(1024)	<=	VN_out_sigd(118);
CN_in_sigd(2480)	<=	VN_out_sigd(118);
CN_in_sigd(2784)	<=	VN_out_sigd(118);
CN_in_sigd(3976)	<=	VN_out_sigd(118);
CN_in_sigd(1032)	<=	VN_out_sigd(119);
CN_in_sigd(2488)	<=	VN_out_sigd(119);
CN_in_sigd(2792)	<=	VN_out_sigd(119);
CN_in_sigd(3984)	<=	VN_out_sigd(119);
CN_in_sigd(1040)	<=	VN_out_sigd(120);
CN_in_sigd(2496)	<=	VN_out_sigd(120);
CN_in_sigd(2800)	<=	VN_out_sigd(120);
CN_in_sigd(3992)	<=	VN_out_sigd(120);
CN_in_sigd(1048)	<=	VN_out_sigd(121);
CN_in_sigd(2504)	<=	VN_out_sigd(121);
CN_in_sigd(2808)	<=	VN_out_sigd(121);
CN_in_sigd(4000)	<=	VN_out_sigd(121);
CN_in_sigd(1056)	<=	VN_out_sigd(122);
CN_in_sigd(2512)	<=	VN_out_sigd(122);
CN_in_sigd(2816)	<=	VN_out_sigd(122);
CN_in_sigd(4008)	<=	VN_out_sigd(122);
CN_in_sigd(1064)	<=	VN_out_sigd(123);
CN_in_sigd(2520)	<=	VN_out_sigd(123);
CN_in_sigd(2824)	<=	VN_out_sigd(123);
CN_in_sigd(4016)	<=	VN_out_sigd(123);
CN_in_sigd(1072)	<=	VN_out_sigd(124);
CN_in_sigd(2528)	<=	VN_out_sigd(124);
CN_in_sigd(2832)	<=	VN_out_sigd(124);
CN_in_sigd(4024)	<=	VN_out_sigd(124);
CN_in_sigd(1080)	<=	VN_out_sigd(125);
CN_in_sigd(2536)	<=	VN_out_sigd(125);
CN_in_sigd(2840)	<=	VN_out_sigd(125);
CN_in_sigd(4032)	<=	VN_out_sigd(125);
CN_in_sigd(1088)	<=	VN_out_sigd(126);
CN_in_sigd(2544)	<=	VN_out_sigd(126);
CN_in_sigd(2848)	<=	VN_out_sigd(126);
CN_in_sigd(4040)	<=	VN_out_sigd(126);
CN_in_sigd(1096)	<=	VN_out_sigd(127);
CN_in_sigd(2552)	<=	VN_out_sigd(127);
CN_in_sigd(2856)	<=	VN_out_sigd(127);
CN_in_sigd(4048)	<=	VN_out_sigd(127);
CN_in_sigd(1104)	<=	VN_out_sigd(128);
CN_in_sigd(2560)	<=	VN_out_sigd(128);
CN_in_sigd(2864)	<=	VN_out_sigd(128);
CN_in_sigd(4056)	<=	VN_out_sigd(128);
CN_in_sigd(1112)	<=	VN_out_sigd(129);
CN_in_sigd(2568)	<=	VN_out_sigd(129);
CN_in_sigd(2872)	<=	VN_out_sigd(129);
CN_in_sigd(4064)	<=	VN_out_sigd(129);
CN_in_sigd(1120)	<=	VN_out_sigd(130);
CN_in_sigd(2576)	<=	VN_out_sigd(130);
CN_in_sigd(2880)	<=	VN_out_sigd(130);
CN_in_sigd(4072)	<=	VN_out_sigd(130);
CN_in_sigd(1128)	<=	VN_out_sigd(131);
CN_in_sigd(2584)	<=	VN_out_sigd(131);
CN_in_sigd(2888)	<=	VN_out_sigd(131);
CN_in_sigd(4080)	<=	VN_out_sigd(131);
CN_in_sigd(1136)	<=	VN_out_sigd(132);
CN_in_sigd(2160)	<=	VN_out_sigd(132);
CN_in_sigd(2896)	<=	VN_out_sigd(132);
CN_in_sigd(4088)	<=	VN_out_sigd(132);
CN_in_sigd(1144)	<=	VN_out_sigd(133);
CN_in_sigd(2168)	<=	VN_out_sigd(133);
CN_in_sigd(2904)	<=	VN_out_sigd(133);
CN_in_sigd(4096)	<=	VN_out_sigd(133);
CN_in_sigd(1152)	<=	VN_out_sigd(134);
CN_in_sigd(2176)	<=	VN_out_sigd(134);
CN_in_sigd(2912)	<=	VN_out_sigd(134);
CN_in_sigd(4104)	<=	VN_out_sigd(134);
CN_in_sigd(1160)	<=	VN_out_sigd(135);
CN_in_sigd(2184)	<=	VN_out_sigd(135);
CN_in_sigd(2920)	<=	VN_out_sigd(135);
CN_in_sigd(4112)	<=	VN_out_sigd(135);
CN_in_sigd(1168)	<=	VN_out_sigd(136);
CN_in_sigd(2192)	<=	VN_out_sigd(136);
CN_in_sigd(2928)	<=	VN_out_sigd(136);
CN_in_sigd(4120)	<=	VN_out_sigd(136);
CN_in_sigd(1176)	<=	VN_out_sigd(137);
CN_in_sigd(2200)	<=	VN_out_sigd(137);
CN_in_sigd(2936)	<=	VN_out_sigd(137);
CN_in_sigd(4128)	<=	VN_out_sigd(137);
CN_in_sigd(1184)	<=	VN_out_sigd(138);
CN_in_sigd(2208)	<=	VN_out_sigd(138);
CN_in_sigd(2944)	<=	VN_out_sigd(138);
CN_in_sigd(4136)	<=	VN_out_sigd(138);
CN_in_sigd(1192)	<=	VN_out_sigd(139);
CN_in_sigd(2216)	<=	VN_out_sigd(139);
CN_in_sigd(2952)	<=	VN_out_sigd(139);
CN_in_sigd(4144)	<=	VN_out_sigd(139);
CN_in_sigd(1200)	<=	VN_out_sigd(140);
CN_in_sigd(2224)	<=	VN_out_sigd(140);
CN_in_sigd(2960)	<=	VN_out_sigd(140);
CN_in_sigd(4152)	<=	VN_out_sigd(140);
CN_in_sigd(1208)	<=	VN_out_sigd(141);
CN_in_sigd(2232)	<=	VN_out_sigd(141);
CN_in_sigd(2968)	<=	VN_out_sigd(141);
CN_in_sigd(4160)	<=	VN_out_sigd(141);
CN_in_sigd(1216)	<=	VN_out_sigd(142);
CN_in_sigd(2240)	<=	VN_out_sigd(142);
CN_in_sigd(2976)	<=	VN_out_sigd(142);
CN_in_sigd(4168)	<=	VN_out_sigd(142);
CN_in_sigd(1224)	<=	VN_out_sigd(143);
CN_in_sigd(2248)	<=	VN_out_sigd(143);
CN_in_sigd(2984)	<=	VN_out_sigd(143);
CN_in_sigd(4176)	<=	VN_out_sigd(143);
CN_in_sigd(1232)	<=	VN_out_sigd(144);
CN_in_sigd(2256)	<=	VN_out_sigd(144);
CN_in_sigd(2992)	<=	VN_out_sigd(144);
CN_in_sigd(4184)	<=	VN_out_sigd(144);
CN_in_sigd(1240)	<=	VN_out_sigd(145);
CN_in_sigd(2264)	<=	VN_out_sigd(145);
CN_in_sigd(3000)	<=	VN_out_sigd(145);
CN_in_sigd(4192)	<=	VN_out_sigd(145);
CN_in_sigd(1248)	<=	VN_out_sigd(146);
CN_in_sigd(2272)	<=	VN_out_sigd(146);
CN_in_sigd(3008)	<=	VN_out_sigd(146);
CN_in_sigd(4200)	<=	VN_out_sigd(146);
CN_in_sigd(1256)	<=	VN_out_sigd(147);
CN_in_sigd(2280)	<=	VN_out_sigd(147);
CN_in_sigd(3016)	<=	VN_out_sigd(147);
CN_in_sigd(4208)	<=	VN_out_sigd(147);
CN_in_sigd(1264)	<=	VN_out_sigd(148);
CN_in_sigd(2288)	<=	VN_out_sigd(148);
CN_in_sigd(2592)	<=	VN_out_sigd(148);
CN_in_sigd(4216)	<=	VN_out_sigd(148);
CN_in_sigd(1272)	<=	VN_out_sigd(149);
CN_in_sigd(2296)	<=	VN_out_sigd(149);
CN_in_sigd(2600)	<=	VN_out_sigd(149);
CN_in_sigd(4224)	<=	VN_out_sigd(149);
CN_in_sigd(1280)	<=	VN_out_sigd(150);
CN_in_sigd(2304)	<=	VN_out_sigd(150);
CN_in_sigd(2608)	<=	VN_out_sigd(150);
CN_in_sigd(4232)	<=	VN_out_sigd(150);
CN_in_sigd(1288)	<=	VN_out_sigd(151);
CN_in_sigd(2312)	<=	VN_out_sigd(151);
CN_in_sigd(2616)	<=	VN_out_sigd(151);
CN_in_sigd(4240)	<=	VN_out_sigd(151);
CN_in_sigd(864)	<=	VN_out_sigd(152);
CN_in_sigd(2320)	<=	VN_out_sigd(152);
CN_in_sigd(2624)	<=	VN_out_sigd(152);
CN_in_sigd(4248)	<=	VN_out_sigd(152);
CN_in_sigd(872)	<=	VN_out_sigd(153);
CN_in_sigd(2328)	<=	VN_out_sigd(153);
CN_in_sigd(2632)	<=	VN_out_sigd(153);
CN_in_sigd(4256)	<=	VN_out_sigd(153);
CN_in_sigd(880)	<=	VN_out_sigd(154);
CN_in_sigd(2336)	<=	VN_out_sigd(154);
CN_in_sigd(2640)	<=	VN_out_sigd(154);
CN_in_sigd(4264)	<=	VN_out_sigd(154);
CN_in_sigd(888)	<=	VN_out_sigd(155);
CN_in_sigd(2344)	<=	VN_out_sigd(155);
CN_in_sigd(2648)	<=	VN_out_sigd(155);
CN_in_sigd(4272)	<=	VN_out_sigd(155);
CN_in_sigd(896)	<=	VN_out_sigd(156);
CN_in_sigd(2352)	<=	VN_out_sigd(156);
CN_in_sigd(2656)	<=	VN_out_sigd(156);
CN_in_sigd(4280)	<=	VN_out_sigd(156);
CN_in_sigd(904)	<=	VN_out_sigd(157);
CN_in_sigd(2360)	<=	VN_out_sigd(157);
CN_in_sigd(2664)	<=	VN_out_sigd(157);
CN_in_sigd(4288)	<=	VN_out_sigd(157);
CN_in_sigd(912)	<=	VN_out_sigd(158);
CN_in_sigd(2368)	<=	VN_out_sigd(158);
CN_in_sigd(2672)	<=	VN_out_sigd(158);
CN_in_sigd(4296)	<=	VN_out_sigd(158);
CN_in_sigd(920)	<=	VN_out_sigd(159);
CN_in_sigd(2376)	<=	VN_out_sigd(159);
CN_in_sigd(2680)	<=	VN_out_sigd(159);
CN_in_sigd(4304)	<=	VN_out_sigd(159);
CN_in_sigd(928)	<=	VN_out_sigd(160);
CN_in_sigd(2384)	<=	VN_out_sigd(160);
CN_in_sigd(2688)	<=	VN_out_sigd(160);
CN_in_sigd(4312)	<=	VN_out_sigd(160);
CN_in_sigd(936)	<=	VN_out_sigd(161);
CN_in_sigd(2392)	<=	VN_out_sigd(161);
CN_in_sigd(2696)	<=	VN_out_sigd(161);
CN_in_sigd(3888)	<=	VN_out_sigd(161);
CN_in_sigd(1265)	<=	VN_out_sigd(162);
CN_in_sigd(1985)	<=	VN_out_sigd(162);
CN_in_sigd(3025)	<=	VN_out_sigd(162);
CN_in_sigd(5049)	<=	VN_out_sigd(162);
CN_in_sigd(1273)	<=	VN_out_sigd(163);
CN_in_sigd(1993)	<=	VN_out_sigd(163);
CN_in_sigd(3033)	<=	VN_out_sigd(163);
CN_in_sigd(5057)	<=	VN_out_sigd(163);
CN_in_sigd(1281)	<=	VN_out_sigd(164);
CN_in_sigd(2001)	<=	VN_out_sigd(164);
CN_in_sigd(3041)	<=	VN_out_sigd(164);
CN_in_sigd(5065)	<=	VN_out_sigd(164);
CN_in_sigd(1289)	<=	VN_out_sigd(165);
CN_in_sigd(2009)	<=	VN_out_sigd(165);
CN_in_sigd(3049)	<=	VN_out_sigd(165);
CN_in_sigd(5073)	<=	VN_out_sigd(165);
CN_in_sigd(865)	<=	VN_out_sigd(166);
CN_in_sigd(2017)	<=	VN_out_sigd(166);
CN_in_sigd(3057)	<=	VN_out_sigd(166);
CN_in_sigd(5081)	<=	VN_out_sigd(166);
CN_in_sigd(873)	<=	VN_out_sigd(167);
CN_in_sigd(2025)	<=	VN_out_sigd(167);
CN_in_sigd(3065)	<=	VN_out_sigd(167);
CN_in_sigd(5089)	<=	VN_out_sigd(167);
CN_in_sigd(881)	<=	VN_out_sigd(168);
CN_in_sigd(2033)	<=	VN_out_sigd(168);
CN_in_sigd(3073)	<=	VN_out_sigd(168);
CN_in_sigd(5097)	<=	VN_out_sigd(168);
CN_in_sigd(889)	<=	VN_out_sigd(169);
CN_in_sigd(2041)	<=	VN_out_sigd(169);
CN_in_sigd(3081)	<=	VN_out_sigd(169);
CN_in_sigd(5105)	<=	VN_out_sigd(169);
CN_in_sigd(897)	<=	VN_out_sigd(170);
CN_in_sigd(2049)	<=	VN_out_sigd(170);
CN_in_sigd(3089)	<=	VN_out_sigd(170);
CN_in_sigd(5113)	<=	VN_out_sigd(170);
CN_in_sigd(905)	<=	VN_out_sigd(171);
CN_in_sigd(2057)	<=	VN_out_sigd(171);
CN_in_sigd(3097)	<=	VN_out_sigd(171);
CN_in_sigd(5121)	<=	VN_out_sigd(171);
CN_in_sigd(913)	<=	VN_out_sigd(172);
CN_in_sigd(2065)	<=	VN_out_sigd(172);
CN_in_sigd(3105)	<=	VN_out_sigd(172);
CN_in_sigd(5129)	<=	VN_out_sigd(172);
CN_in_sigd(921)	<=	VN_out_sigd(173);
CN_in_sigd(2073)	<=	VN_out_sigd(173);
CN_in_sigd(3113)	<=	VN_out_sigd(173);
CN_in_sigd(5137)	<=	VN_out_sigd(173);
CN_in_sigd(929)	<=	VN_out_sigd(174);
CN_in_sigd(2081)	<=	VN_out_sigd(174);
CN_in_sigd(3121)	<=	VN_out_sigd(174);
CN_in_sigd(5145)	<=	VN_out_sigd(174);
CN_in_sigd(937)	<=	VN_out_sigd(175);
CN_in_sigd(2089)	<=	VN_out_sigd(175);
CN_in_sigd(3129)	<=	VN_out_sigd(175);
CN_in_sigd(5153)	<=	VN_out_sigd(175);
CN_in_sigd(945)	<=	VN_out_sigd(176);
CN_in_sigd(2097)	<=	VN_out_sigd(176);
CN_in_sigd(3137)	<=	VN_out_sigd(176);
CN_in_sigd(5161)	<=	VN_out_sigd(176);
CN_in_sigd(953)	<=	VN_out_sigd(177);
CN_in_sigd(2105)	<=	VN_out_sigd(177);
CN_in_sigd(3145)	<=	VN_out_sigd(177);
CN_in_sigd(5169)	<=	VN_out_sigd(177);
CN_in_sigd(961)	<=	VN_out_sigd(178);
CN_in_sigd(2113)	<=	VN_out_sigd(178);
CN_in_sigd(3153)	<=	VN_out_sigd(178);
CN_in_sigd(5177)	<=	VN_out_sigd(178);
CN_in_sigd(969)	<=	VN_out_sigd(179);
CN_in_sigd(2121)	<=	VN_out_sigd(179);
CN_in_sigd(3161)	<=	VN_out_sigd(179);
CN_in_sigd(4753)	<=	VN_out_sigd(179);
CN_in_sigd(977)	<=	VN_out_sigd(180);
CN_in_sigd(2129)	<=	VN_out_sigd(180);
CN_in_sigd(3169)	<=	VN_out_sigd(180);
CN_in_sigd(4761)	<=	VN_out_sigd(180);
CN_in_sigd(985)	<=	VN_out_sigd(181);
CN_in_sigd(2137)	<=	VN_out_sigd(181);
CN_in_sigd(3177)	<=	VN_out_sigd(181);
CN_in_sigd(4769)	<=	VN_out_sigd(181);
CN_in_sigd(993)	<=	VN_out_sigd(182);
CN_in_sigd(2145)	<=	VN_out_sigd(182);
CN_in_sigd(3185)	<=	VN_out_sigd(182);
CN_in_sigd(4777)	<=	VN_out_sigd(182);
CN_in_sigd(1001)	<=	VN_out_sigd(183);
CN_in_sigd(2153)	<=	VN_out_sigd(183);
CN_in_sigd(3193)	<=	VN_out_sigd(183);
CN_in_sigd(4785)	<=	VN_out_sigd(183);
CN_in_sigd(1009)	<=	VN_out_sigd(184);
CN_in_sigd(1729)	<=	VN_out_sigd(184);
CN_in_sigd(3201)	<=	VN_out_sigd(184);
CN_in_sigd(4793)	<=	VN_out_sigd(184);
CN_in_sigd(1017)	<=	VN_out_sigd(185);
CN_in_sigd(1737)	<=	VN_out_sigd(185);
CN_in_sigd(3209)	<=	VN_out_sigd(185);
CN_in_sigd(4801)	<=	VN_out_sigd(185);
CN_in_sigd(1025)	<=	VN_out_sigd(186);
CN_in_sigd(1745)	<=	VN_out_sigd(186);
CN_in_sigd(3217)	<=	VN_out_sigd(186);
CN_in_sigd(4809)	<=	VN_out_sigd(186);
CN_in_sigd(1033)	<=	VN_out_sigd(187);
CN_in_sigd(1753)	<=	VN_out_sigd(187);
CN_in_sigd(3225)	<=	VN_out_sigd(187);
CN_in_sigd(4817)	<=	VN_out_sigd(187);
CN_in_sigd(1041)	<=	VN_out_sigd(188);
CN_in_sigd(1761)	<=	VN_out_sigd(188);
CN_in_sigd(3233)	<=	VN_out_sigd(188);
CN_in_sigd(4825)	<=	VN_out_sigd(188);
CN_in_sigd(1049)	<=	VN_out_sigd(189);
CN_in_sigd(1769)	<=	VN_out_sigd(189);
CN_in_sigd(3241)	<=	VN_out_sigd(189);
CN_in_sigd(4833)	<=	VN_out_sigd(189);
CN_in_sigd(1057)	<=	VN_out_sigd(190);
CN_in_sigd(1777)	<=	VN_out_sigd(190);
CN_in_sigd(3249)	<=	VN_out_sigd(190);
CN_in_sigd(4841)	<=	VN_out_sigd(190);
CN_in_sigd(1065)	<=	VN_out_sigd(191);
CN_in_sigd(1785)	<=	VN_out_sigd(191);
CN_in_sigd(3257)	<=	VN_out_sigd(191);
CN_in_sigd(4849)	<=	VN_out_sigd(191);
CN_in_sigd(1073)	<=	VN_out_sigd(192);
CN_in_sigd(1793)	<=	VN_out_sigd(192);
CN_in_sigd(3265)	<=	VN_out_sigd(192);
CN_in_sigd(4857)	<=	VN_out_sigd(192);
CN_in_sigd(1081)	<=	VN_out_sigd(193);
CN_in_sigd(1801)	<=	VN_out_sigd(193);
CN_in_sigd(3273)	<=	VN_out_sigd(193);
CN_in_sigd(4865)	<=	VN_out_sigd(193);
CN_in_sigd(1089)	<=	VN_out_sigd(194);
CN_in_sigd(1809)	<=	VN_out_sigd(194);
CN_in_sigd(3281)	<=	VN_out_sigd(194);
CN_in_sigd(4873)	<=	VN_out_sigd(194);
CN_in_sigd(1097)	<=	VN_out_sigd(195);
CN_in_sigd(1817)	<=	VN_out_sigd(195);
CN_in_sigd(3289)	<=	VN_out_sigd(195);
CN_in_sigd(4881)	<=	VN_out_sigd(195);
CN_in_sigd(1105)	<=	VN_out_sigd(196);
CN_in_sigd(1825)	<=	VN_out_sigd(196);
CN_in_sigd(3297)	<=	VN_out_sigd(196);
CN_in_sigd(4889)	<=	VN_out_sigd(196);
CN_in_sigd(1113)	<=	VN_out_sigd(197);
CN_in_sigd(1833)	<=	VN_out_sigd(197);
CN_in_sigd(3305)	<=	VN_out_sigd(197);
CN_in_sigd(4897)	<=	VN_out_sigd(197);
CN_in_sigd(1121)	<=	VN_out_sigd(198);
CN_in_sigd(1841)	<=	VN_out_sigd(198);
CN_in_sigd(3313)	<=	VN_out_sigd(198);
CN_in_sigd(4905)	<=	VN_out_sigd(198);
CN_in_sigd(1129)	<=	VN_out_sigd(199);
CN_in_sigd(1849)	<=	VN_out_sigd(199);
CN_in_sigd(3321)	<=	VN_out_sigd(199);
CN_in_sigd(4913)	<=	VN_out_sigd(199);
CN_in_sigd(1137)	<=	VN_out_sigd(200);
CN_in_sigd(1857)	<=	VN_out_sigd(200);
CN_in_sigd(3329)	<=	VN_out_sigd(200);
CN_in_sigd(4921)	<=	VN_out_sigd(200);
CN_in_sigd(1145)	<=	VN_out_sigd(201);
CN_in_sigd(1865)	<=	VN_out_sigd(201);
CN_in_sigd(3337)	<=	VN_out_sigd(201);
CN_in_sigd(4929)	<=	VN_out_sigd(201);
CN_in_sigd(1153)	<=	VN_out_sigd(202);
CN_in_sigd(1873)	<=	VN_out_sigd(202);
CN_in_sigd(3345)	<=	VN_out_sigd(202);
CN_in_sigd(4937)	<=	VN_out_sigd(202);
CN_in_sigd(1161)	<=	VN_out_sigd(203);
CN_in_sigd(1881)	<=	VN_out_sigd(203);
CN_in_sigd(3353)	<=	VN_out_sigd(203);
CN_in_sigd(4945)	<=	VN_out_sigd(203);
CN_in_sigd(1169)	<=	VN_out_sigd(204);
CN_in_sigd(1889)	<=	VN_out_sigd(204);
CN_in_sigd(3361)	<=	VN_out_sigd(204);
CN_in_sigd(4953)	<=	VN_out_sigd(204);
CN_in_sigd(1177)	<=	VN_out_sigd(205);
CN_in_sigd(1897)	<=	VN_out_sigd(205);
CN_in_sigd(3369)	<=	VN_out_sigd(205);
CN_in_sigd(4961)	<=	VN_out_sigd(205);
CN_in_sigd(1185)	<=	VN_out_sigd(206);
CN_in_sigd(1905)	<=	VN_out_sigd(206);
CN_in_sigd(3377)	<=	VN_out_sigd(206);
CN_in_sigd(4969)	<=	VN_out_sigd(206);
CN_in_sigd(1193)	<=	VN_out_sigd(207);
CN_in_sigd(1913)	<=	VN_out_sigd(207);
CN_in_sigd(3385)	<=	VN_out_sigd(207);
CN_in_sigd(4977)	<=	VN_out_sigd(207);
CN_in_sigd(1201)	<=	VN_out_sigd(208);
CN_in_sigd(1921)	<=	VN_out_sigd(208);
CN_in_sigd(3393)	<=	VN_out_sigd(208);
CN_in_sigd(4985)	<=	VN_out_sigd(208);
CN_in_sigd(1209)	<=	VN_out_sigd(209);
CN_in_sigd(1929)	<=	VN_out_sigd(209);
CN_in_sigd(3401)	<=	VN_out_sigd(209);
CN_in_sigd(4993)	<=	VN_out_sigd(209);
CN_in_sigd(1217)	<=	VN_out_sigd(210);
CN_in_sigd(1937)	<=	VN_out_sigd(210);
CN_in_sigd(3409)	<=	VN_out_sigd(210);
CN_in_sigd(5001)	<=	VN_out_sigd(210);
CN_in_sigd(1225)	<=	VN_out_sigd(211);
CN_in_sigd(1945)	<=	VN_out_sigd(211);
CN_in_sigd(3417)	<=	VN_out_sigd(211);
CN_in_sigd(5009)	<=	VN_out_sigd(211);
CN_in_sigd(1233)	<=	VN_out_sigd(212);
CN_in_sigd(1953)	<=	VN_out_sigd(212);
CN_in_sigd(3425)	<=	VN_out_sigd(212);
CN_in_sigd(5017)	<=	VN_out_sigd(212);
CN_in_sigd(1241)	<=	VN_out_sigd(213);
CN_in_sigd(1961)	<=	VN_out_sigd(213);
CN_in_sigd(3433)	<=	VN_out_sigd(213);
CN_in_sigd(5025)	<=	VN_out_sigd(213);
CN_in_sigd(1249)	<=	VN_out_sigd(214);
CN_in_sigd(1969)	<=	VN_out_sigd(214);
CN_in_sigd(3441)	<=	VN_out_sigd(214);
CN_in_sigd(5033)	<=	VN_out_sigd(214);
CN_in_sigd(1257)	<=	VN_out_sigd(215);
CN_in_sigd(1977)	<=	VN_out_sigd(215);
CN_in_sigd(3449)	<=	VN_out_sigd(215);
CN_in_sigd(5041)	<=	VN_out_sigd(215);
CN_in_sigd(217)	<=	VN_out_sigd(216);
CN_in_sigd(1457)	<=	VN_out_sigd(216);
CN_in_sigd(3833)	<=	VN_out_sigd(216);
CN_in_sigd(4721)	<=	VN_out_sigd(216);
CN_in_sigd(225)	<=	VN_out_sigd(217);
CN_in_sigd(1465)	<=	VN_out_sigd(217);
CN_in_sigd(3841)	<=	VN_out_sigd(217);
CN_in_sigd(4729)	<=	VN_out_sigd(217);
CN_in_sigd(233)	<=	VN_out_sigd(218);
CN_in_sigd(1473)	<=	VN_out_sigd(218);
CN_in_sigd(3849)	<=	VN_out_sigd(218);
CN_in_sigd(4737)	<=	VN_out_sigd(218);
CN_in_sigd(241)	<=	VN_out_sigd(219);
CN_in_sigd(1481)	<=	VN_out_sigd(219);
CN_in_sigd(3857)	<=	VN_out_sigd(219);
CN_in_sigd(4745)	<=	VN_out_sigd(219);
CN_in_sigd(249)	<=	VN_out_sigd(220);
CN_in_sigd(1489)	<=	VN_out_sigd(220);
CN_in_sigd(3865)	<=	VN_out_sigd(220);
CN_in_sigd(4321)	<=	VN_out_sigd(220);
CN_in_sigd(257)	<=	VN_out_sigd(221);
CN_in_sigd(1497)	<=	VN_out_sigd(221);
CN_in_sigd(3873)	<=	VN_out_sigd(221);
CN_in_sigd(4329)	<=	VN_out_sigd(221);
CN_in_sigd(265)	<=	VN_out_sigd(222);
CN_in_sigd(1505)	<=	VN_out_sigd(222);
CN_in_sigd(3881)	<=	VN_out_sigd(222);
CN_in_sigd(4337)	<=	VN_out_sigd(222);
CN_in_sigd(273)	<=	VN_out_sigd(223);
CN_in_sigd(1513)	<=	VN_out_sigd(223);
CN_in_sigd(3457)	<=	VN_out_sigd(223);
CN_in_sigd(4345)	<=	VN_out_sigd(223);
CN_in_sigd(281)	<=	VN_out_sigd(224);
CN_in_sigd(1521)	<=	VN_out_sigd(224);
CN_in_sigd(3465)	<=	VN_out_sigd(224);
CN_in_sigd(4353)	<=	VN_out_sigd(224);
CN_in_sigd(289)	<=	VN_out_sigd(225);
CN_in_sigd(1529)	<=	VN_out_sigd(225);
CN_in_sigd(3473)	<=	VN_out_sigd(225);
CN_in_sigd(4361)	<=	VN_out_sigd(225);
CN_in_sigd(297)	<=	VN_out_sigd(226);
CN_in_sigd(1537)	<=	VN_out_sigd(226);
CN_in_sigd(3481)	<=	VN_out_sigd(226);
CN_in_sigd(4369)	<=	VN_out_sigd(226);
CN_in_sigd(305)	<=	VN_out_sigd(227);
CN_in_sigd(1545)	<=	VN_out_sigd(227);
CN_in_sigd(3489)	<=	VN_out_sigd(227);
CN_in_sigd(4377)	<=	VN_out_sigd(227);
CN_in_sigd(313)	<=	VN_out_sigd(228);
CN_in_sigd(1553)	<=	VN_out_sigd(228);
CN_in_sigd(3497)	<=	VN_out_sigd(228);
CN_in_sigd(4385)	<=	VN_out_sigd(228);
CN_in_sigd(321)	<=	VN_out_sigd(229);
CN_in_sigd(1561)	<=	VN_out_sigd(229);
CN_in_sigd(3505)	<=	VN_out_sigd(229);
CN_in_sigd(4393)	<=	VN_out_sigd(229);
CN_in_sigd(329)	<=	VN_out_sigd(230);
CN_in_sigd(1569)	<=	VN_out_sigd(230);
CN_in_sigd(3513)	<=	VN_out_sigd(230);
CN_in_sigd(4401)	<=	VN_out_sigd(230);
CN_in_sigd(337)	<=	VN_out_sigd(231);
CN_in_sigd(1577)	<=	VN_out_sigd(231);
CN_in_sigd(3521)	<=	VN_out_sigd(231);
CN_in_sigd(4409)	<=	VN_out_sigd(231);
CN_in_sigd(345)	<=	VN_out_sigd(232);
CN_in_sigd(1585)	<=	VN_out_sigd(232);
CN_in_sigd(3529)	<=	VN_out_sigd(232);
CN_in_sigd(4417)	<=	VN_out_sigd(232);
CN_in_sigd(353)	<=	VN_out_sigd(233);
CN_in_sigd(1593)	<=	VN_out_sigd(233);
CN_in_sigd(3537)	<=	VN_out_sigd(233);
CN_in_sigd(4425)	<=	VN_out_sigd(233);
CN_in_sigd(361)	<=	VN_out_sigd(234);
CN_in_sigd(1601)	<=	VN_out_sigd(234);
CN_in_sigd(3545)	<=	VN_out_sigd(234);
CN_in_sigd(4433)	<=	VN_out_sigd(234);
CN_in_sigd(369)	<=	VN_out_sigd(235);
CN_in_sigd(1609)	<=	VN_out_sigd(235);
CN_in_sigd(3553)	<=	VN_out_sigd(235);
CN_in_sigd(4441)	<=	VN_out_sigd(235);
CN_in_sigd(377)	<=	VN_out_sigd(236);
CN_in_sigd(1617)	<=	VN_out_sigd(236);
CN_in_sigd(3561)	<=	VN_out_sigd(236);
CN_in_sigd(4449)	<=	VN_out_sigd(236);
CN_in_sigd(385)	<=	VN_out_sigd(237);
CN_in_sigd(1625)	<=	VN_out_sigd(237);
CN_in_sigd(3569)	<=	VN_out_sigd(237);
CN_in_sigd(4457)	<=	VN_out_sigd(237);
CN_in_sigd(393)	<=	VN_out_sigd(238);
CN_in_sigd(1633)	<=	VN_out_sigd(238);
CN_in_sigd(3577)	<=	VN_out_sigd(238);
CN_in_sigd(4465)	<=	VN_out_sigd(238);
CN_in_sigd(401)	<=	VN_out_sigd(239);
CN_in_sigd(1641)	<=	VN_out_sigd(239);
CN_in_sigd(3585)	<=	VN_out_sigd(239);
CN_in_sigd(4473)	<=	VN_out_sigd(239);
CN_in_sigd(409)	<=	VN_out_sigd(240);
CN_in_sigd(1649)	<=	VN_out_sigd(240);
CN_in_sigd(3593)	<=	VN_out_sigd(240);
CN_in_sigd(4481)	<=	VN_out_sigd(240);
CN_in_sigd(417)	<=	VN_out_sigd(241);
CN_in_sigd(1657)	<=	VN_out_sigd(241);
CN_in_sigd(3601)	<=	VN_out_sigd(241);
CN_in_sigd(4489)	<=	VN_out_sigd(241);
CN_in_sigd(425)	<=	VN_out_sigd(242);
CN_in_sigd(1665)	<=	VN_out_sigd(242);
CN_in_sigd(3609)	<=	VN_out_sigd(242);
CN_in_sigd(4497)	<=	VN_out_sigd(242);
CN_in_sigd(1)	<=	VN_out_sigd(243);
CN_in_sigd(1673)	<=	VN_out_sigd(243);
CN_in_sigd(3617)	<=	VN_out_sigd(243);
CN_in_sigd(4505)	<=	VN_out_sigd(243);
CN_in_sigd(9)	<=	VN_out_sigd(244);
CN_in_sigd(1681)	<=	VN_out_sigd(244);
CN_in_sigd(3625)	<=	VN_out_sigd(244);
CN_in_sigd(4513)	<=	VN_out_sigd(244);
CN_in_sigd(17)	<=	VN_out_sigd(245);
CN_in_sigd(1689)	<=	VN_out_sigd(245);
CN_in_sigd(3633)	<=	VN_out_sigd(245);
CN_in_sigd(4521)	<=	VN_out_sigd(245);
CN_in_sigd(25)	<=	VN_out_sigd(246);
CN_in_sigd(1697)	<=	VN_out_sigd(246);
CN_in_sigd(3641)	<=	VN_out_sigd(246);
CN_in_sigd(4529)	<=	VN_out_sigd(246);
CN_in_sigd(33)	<=	VN_out_sigd(247);
CN_in_sigd(1705)	<=	VN_out_sigd(247);
CN_in_sigd(3649)	<=	VN_out_sigd(247);
CN_in_sigd(4537)	<=	VN_out_sigd(247);
CN_in_sigd(41)	<=	VN_out_sigd(248);
CN_in_sigd(1713)	<=	VN_out_sigd(248);
CN_in_sigd(3657)	<=	VN_out_sigd(248);
CN_in_sigd(4545)	<=	VN_out_sigd(248);
CN_in_sigd(49)	<=	VN_out_sigd(249);
CN_in_sigd(1721)	<=	VN_out_sigd(249);
CN_in_sigd(3665)	<=	VN_out_sigd(249);
CN_in_sigd(4553)	<=	VN_out_sigd(249);
CN_in_sigd(57)	<=	VN_out_sigd(250);
CN_in_sigd(1297)	<=	VN_out_sigd(250);
CN_in_sigd(3673)	<=	VN_out_sigd(250);
CN_in_sigd(4561)	<=	VN_out_sigd(250);
CN_in_sigd(65)	<=	VN_out_sigd(251);
CN_in_sigd(1305)	<=	VN_out_sigd(251);
CN_in_sigd(3681)	<=	VN_out_sigd(251);
CN_in_sigd(4569)	<=	VN_out_sigd(251);
CN_in_sigd(73)	<=	VN_out_sigd(252);
CN_in_sigd(1313)	<=	VN_out_sigd(252);
CN_in_sigd(3689)	<=	VN_out_sigd(252);
CN_in_sigd(4577)	<=	VN_out_sigd(252);
CN_in_sigd(81)	<=	VN_out_sigd(253);
CN_in_sigd(1321)	<=	VN_out_sigd(253);
CN_in_sigd(3697)	<=	VN_out_sigd(253);
CN_in_sigd(4585)	<=	VN_out_sigd(253);
CN_in_sigd(89)	<=	VN_out_sigd(254);
CN_in_sigd(1329)	<=	VN_out_sigd(254);
CN_in_sigd(3705)	<=	VN_out_sigd(254);
CN_in_sigd(4593)	<=	VN_out_sigd(254);
CN_in_sigd(97)	<=	VN_out_sigd(255);
CN_in_sigd(1337)	<=	VN_out_sigd(255);
CN_in_sigd(3713)	<=	VN_out_sigd(255);
CN_in_sigd(4601)	<=	VN_out_sigd(255);
CN_in_sigd(105)	<=	VN_out_sigd(256);
CN_in_sigd(1345)	<=	VN_out_sigd(256);
CN_in_sigd(3721)	<=	VN_out_sigd(256);
CN_in_sigd(4609)	<=	VN_out_sigd(256);
CN_in_sigd(113)	<=	VN_out_sigd(257);
CN_in_sigd(1353)	<=	VN_out_sigd(257);
CN_in_sigd(3729)	<=	VN_out_sigd(257);
CN_in_sigd(4617)	<=	VN_out_sigd(257);
CN_in_sigd(121)	<=	VN_out_sigd(258);
CN_in_sigd(1361)	<=	VN_out_sigd(258);
CN_in_sigd(3737)	<=	VN_out_sigd(258);
CN_in_sigd(4625)	<=	VN_out_sigd(258);
CN_in_sigd(129)	<=	VN_out_sigd(259);
CN_in_sigd(1369)	<=	VN_out_sigd(259);
CN_in_sigd(3745)	<=	VN_out_sigd(259);
CN_in_sigd(4633)	<=	VN_out_sigd(259);
CN_in_sigd(137)	<=	VN_out_sigd(260);
CN_in_sigd(1377)	<=	VN_out_sigd(260);
CN_in_sigd(3753)	<=	VN_out_sigd(260);
CN_in_sigd(4641)	<=	VN_out_sigd(260);
CN_in_sigd(145)	<=	VN_out_sigd(261);
CN_in_sigd(1385)	<=	VN_out_sigd(261);
CN_in_sigd(3761)	<=	VN_out_sigd(261);
CN_in_sigd(4649)	<=	VN_out_sigd(261);
CN_in_sigd(153)	<=	VN_out_sigd(262);
CN_in_sigd(1393)	<=	VN_out_sigd(262);
CN_in_sigd(3769)	<=	VN_out_sigd(262);
CN_in_sigd(4657)	<=	VN_out_sigd(262);
CN_in_sigd(161)	<=	VN_out_sigd(263);
CN_in_sigd(1401)	<=	VN_out_sigd(263);
CN_in_sigd(3777)	<=	VN_out_sigd(263);
CN_in_sigd(4665)	<=	VN_out_sigd(263);
CN_in_sigd(169)	<=	VN_out_sigd(264);
CN_in_sigd(1409)	<=	VN_out_sigd(264);
CN_in_sigd(3785)	<=	VN_out_sigd(264);
CN_in_sigd(4673)	<=	VN_out_sigd(264);
CN_in_sigd(177)	<=	VN_out_sigd(265);
CN_in_sigd(1417)	<=	VN_out_sigd(265);
CN_in_sigd(3793)	<=	VN_out_sigd(265);
CN_in_sigd(4681)	<=	VN_out_sigd(265);
CN_in_sigd(185)	<=	VN_out_sigd(266);
CN_in_sigd(1425)	<=	VN_out_sigd(266);
CN_in_sigd(3801)	<=	VN_out_sigd(266);
CN_in_sigd(4689)	<=	VN_out_sigd(266);
CN_in_sigd(193)	<=	VN_out_sigd(267);
CN_in_sigd(1433)	<=	VN_out_sigd(267);
CN_in_sigd(3809)	<=	VN_out_sigd(267);
CN_in_sigd(4697)	<=	VN_out_sigd(267);
CN_in_sigd(201)	<=	VN_out_sigd(268);
CN_in_sigd(1441)	<=	VN_out_sigd(268);
CN_in_sigd(3817)	<=	VN_out_sigd(268);
CN_in_sigd(4705)	<=	VN_out_sigd(268);
CN_in_sigd(209)	<=	VN_out_sigd(269);
CN_in_sigd(1449)	<=	VN_out_sigd(269);
CN_in_sigd(3825)	<=	VN_out_sigd(269);
CN_in_sigd(4713)	<=	VN_out_sigd(269);
CN_in_sigd(617)	<=	VN_out_sigd(270);
CN_in_sigd(2513)	<=	VN_out_sigd(270);
CN_in_sigd(2745)	<=	VN_out_sigd(270);
CN_in_sigd(4297)	<=	VN_out_sigd(270);
CN_in_sigd(625)	<=	VN_out_sigd(271);
CN_in_sigd(2521)	<=	VN_out_sigd(271);
CN_in_sigd(2753)	<=	VN_out_sigd(271);
CN_in_sigd(4305)	<=	VN_out_sigd(271);
CN_in_sigd(633)	<=	VN_out_sigd(272);
CN_in_sigd(2529)	<=	VN_out_sigd(272);
CN_in_sigd(2761)	<=	VN_out_sigd(272);
CN_in_sigd(4313)	<=	VN_out_sigd(272);
CN_in_sigd(641)	<=	VN_out_sigd(273);
CN_in_sigd(2537)	<=	VN_out_sigd(273);
CN_in_sigd(2769)	<=	VN_out_sigd(273);
CN_in_sigd(3889)	<=	VN_out_sigd(273);
CN_in_sigd(649)	<=	VN_out_sigd(274);
CN_in_sigd(2545)	<=	VN_out_sigd(274);
CN_in_sigd(2777)	<=	VN_out_sigd(274);
CN_in_sigd(3897)	<=	VN_out_sigd(274);
CN_in_sigd(657)	<=	VN_out_sigd(275);
CN_in_sigd(2553)	<=	VN_out_sigd(275);
CN_in_sigd(2785)	<=	VN_out_sigd(275);
CN_in_sigd(3905)	<=	VN_out_sigd(275);
CN_in_sigd(665)	<=	VN_out_sigd(276);
CN_in_sigd(2561)	<=	VN_out_sigd(276);
CN_in_sigd(2793)	<=	VN_out_sigd(276);
CN_in_sigd(3913)	<=	VN_out_sigd(276);
CN_in_sigd(673)	<=	VN_out_sigd(277);
CN_in_sigd(2569)	<=	VN_out_sigd(277);
CN_in_sigd(2801)	<=	VN_out_sigd(277);
CN_in_sigd(3921)	<=	VN_out_sigd(277);
CN_in_sigd(681)	<=	VN_out_sigd(278);
CN_in_sigd(2577)	<=	VN_out_sigd(278);
CN_in_sigd(2809)	<=	VN_out_sigd(278);
CN_in_sigd(3929)	<=	VN_out_sigd(278);
CN_in_sigd(689)	<=	VN_out_sigd(279);
CN_in_sigd(2585)	<=	VN_out_sigd(279);
CN_in_sigd(2817)	<=	VN_out_sigd(279);
CN_in_sigd(3937)	<=	VN_out_sigd(279);
CN_in_sigd(697)	<=	VN_out_sigd(280);
CN_in_sigd(2161)	<=	VN_out_sigd(280);
CN_in_sigd(2825)	<=	VN_out_sigd(280);
CN_in_sigd(3945)	<=	VN_out_sigd(280);
CN_in_sigd(705)	<=	VN_out_sigd(281);
CN_in_sigd(2169)	<=	VN_out_sigd(281);
CN_in_sigd(2833)	<=	VN_out_sigd(281);
CN_in_sigd(3953)	<=	VN_out_sigd(281);
CN_in_sigd(713)	<=	VN_out_sigd(282);
CN_in_sigd(2177)	<=	VN_out_sigd(282);
CN_in_sigd(2841)	<=	VN_out_sigd(282);
CN_in_sigd(3961)	<=	VN_out_sigd(282);
CN_in_sigd(721)	<=	VN_out_sigd(283);
CN_in_sigd(2185)	<=	VN_out_sigd(283);
CN_in_sigd(2849)	<=	VN_out_sigd(283);
CN_in_sigd(3969)	<=	VN_out_sigd(283);
CN_in_sigd(729)	<=	VN_out_sigd(284);
CN_in_sigd(2193)	<=	VN_out_sigd(284);
CN_in_sigd(2857)	<=	VN_out_sigd(284);
CN_in_sigd(3977)	<=	VN_out_sigd(284);
CN_in_sigd(737)	<=	VN_out_sigd(285);
CN_in_sigd(2201)	<=	VN_out_sigd(285);
CN_in_sigd(2865)	<=	VN_out_sigd(285);
CN_in_sigd(3985)	<=	VN_out_sigd(285);
CN_in_sigd(745)	<=	VN_out_sigd(286);
CN_in_sigd(2209)	<=	VN_out_sigd(286);
CN_in_sigd(2873)	<=	VN_out_sigd(286);
CN_in_sigd(3993)	<=	VN_out_sigd(286);
CN_in_sigd(753)	<=	VN_out_sigd(287);
CN_in_sigd(2217)	<=	VN_out_sigd(287);
CN_in_sigd(2881)	<=	VN_out_sigd(287);
CN_in_sigd(4001)	<=	VN_out_sigd(287);
CN_in_sigd(761)	<=	VN_out_sigd(288);
CN_in_sigd(2225)	<=	VN_out_sigd(288);
CN_in_sigd(2889)	<=	VN_out_sigd(288);
CN_in_sigd(4009)	<=	VN_out_sigd(288);
CN_in_sigd(769)	<=	VN_out_sigd(289);
CN_in_sigd(2233)	<=	VN_out_sigd(289);
CN_in_sigd(2897)	<=	VN_out_sigd(289);
CN_in_sigd(4017)	<=	VN_out_sigd(289);
CN_in_sigd(777)	<=	VN_out_sigd(290);
CN_in_sigd(2241)	<=	VN_out_sigd(290);
CN_in_sigd(2905)	<=	VN_out_sigd(290);
CN_in_sigd(4025)	<=	VN_out_sigd(290);
CN_in_sigd(785)	<=	VN_out_sigd(291);
CN_in_sigd(2249)	<=	VN_out_sigd(291);
CN_in_sigd(2913)	<=	VN_out_sigd(291);
CN_in_sigd(4033)	<=	VN_out_sigd(291);
CN_in_sigd(793)	<=	VN_out_sigd(292);
CN_in_sigd(2257)	<=	VN_out_sigd(292);
CN_in_sigd(2921)	<=	VN_out_sigd(292);
CN_in_sigd(4041)	<=	VN_out_sigd(292);
CN_in_sigd(801)	<=	VN_out_sigd(293);
CN_in_sigd(2265)	<=	VN_out_sigd(293);
CN_in_sigd(2929)	<=	VN_out_sigd(293);
CN_in_sigd(4049)	<=	VN_out_sigd(293);
CN_in_sigd(809)	<=	VN_out_sigd(294);
CN_in_sigd(2273)	<=	VN_out_sigd(294);
CN_in_sigd(2937)	<=	VN_out_sigd(294);
CN_in_sigd(4057)	<=	VN_out_sigd(294);
CN_in_sigd(817)	<=	VN_out_sigd(295);
CN_in_sigd(2281)	<=	VN_out_sigd(295);
CN_in_sigd(2945)	<=	VN_out_sigd(295);
CN_in_sigd(4065)	<=	VN_out_sigd(295);
CN_in_sigd(825)	<=	VN_out_sigd(296);
CN_in_sigd(2289)	<=	VN_out_sigd(296);
CN_in_sigd(2953)	<=	VN_out_sigd(296);
CN_in_sigd(4073)	<=	VN_out_sigd(296);
CN_in_sigd(833)	<=	VN_out_sigd(297);
CN_in_sigd(2297)	<=	VN_out_sigd(297);
CN_in_sigd(2961)	<=	VN_out_sigd(297);
CN_in_sigd(4081)	<=	VN_out_sigd(297);
CN_in_sigd(841)	<=	VN_out_sigd(298);
CN_in_sigd(2305)	<=	VN_out_sigd(298);
CN_in_sigd(2969)	<=	VN_out_sigd(298);
CN_in_sigd(4089)	<=	VN_out_sigd(298);
CN_in_sigd(849)	<=	VN_out_sigd(299);
CN_in_sigd(2313)	<=	VN_out_sigd(299);
CN_in_sigd(2977)	<=	VN_out_sigd(299);
CN_in_sigd(4097)	<=	VN_out_sigd(299);
CN_in_sigd(857)	<=	VN_out_sigd(300);
CN_in_sigd(2321)	<=	VN_out_sigd(300);
CN_in_sigd(2985)	<=	VN_out_sigd(300);
CN_in_sigd(4105)	<=	VN_out_sigd(300);
CN_in_sigd(433)	<=	VN_out_sigd(301);
CN_in_sigd(2329)	<=	VN_out_sigd(301);
CN_in_sigd(2993)	<=	VN_out_sigd(301);
CN_in_sigd(4113)	<=	VN_out_sigd(301);
CN_in_sigd(441)	<=	VN_out_sigd(302);
CN_in_sigd(2337)	<=	VN_out_sigd(302);
CN_in_sigd(3001)	<=	VN_out_sigd(302);
CN_in_sigd(4121)	<=	VN_out_sigd(302);
CN_in_sigd(449)	<=	VN_out_sigd(303);
CN_in_sigd(2345)	<=	VN_out_sigd(303);
CN_in_sigd(3009)	<=	VN_out_sigd(303);
CN_in_sigd(4129)	<=	VN_out_sigd(303);
CN_in_sigd(457)	<=	VN_out_sigd(304);
CN_in_sigd(2353)	<=	VN_out_sigd(304);
CN_in_sigd(3017)	<=	VN_out_sigd(304);
CN_in_sigd(4137)	<=	VN_out_sigd(304);
CN_in_sigd(465)	<=	VN_out_sigd(305);
CN_in_sigd(2361)	<=	VN_out_sigd(305);
CN_in_sigd(2593)	<=	VN_out_sigd(305);
CN_in_sigd(4145)	<=	VN_out_sigd(305);
CN_in_sigd(473)	<=	VN_out_sigd(306);
CN_in_sigd(2369)	<=	VN_out_sigd(306);
CN_in_sigd(2601)	<=	VN_out_sigd(306);
CN_in_sigd(4153)	<=	VN_out_sigd(306);
CN_in_sigd(481)	<=	VN_out_sigd(307);
CN_in_sigd(2377)	<=	VN_out_sigd(307);
CN_in_sigd(2609)	<=	VN_out_sigd(307);
CN_in_sigd(4161)	<=	VN_out_sigd(307);
CN_in_sigd(489)	<=	VN_out_sigd(308);
CN_in_sigd(2385)	<=	VN_out_sigd(308);
CN_in_sigd(2617)	<=	VN_out_sigd(308);
CN_in_sigd(4169)	<=	VN_out_sigd(308);
CN_in_sigd(497)	<=	VN_out_sigd(309);
CN_in_sigd(2393)	<=	VN_out_sigd(309);
CN_in_sigd(2625)	<=	VN_out_sigd(309);
CN_in_sigd(4177)	<=	VN_out_sigd(309);
CN_in_sigd(505)	<=	VN_out_sigd(310);
CN_in_sigd(2401)	<=	VN_out_sigd(310);
CN_in_sigd(2633)	<=	VN_out_sigd(310);
CN_in_sigd(4185)	<=	VN_out_sigd(310);
CN_in_sigd(513)	<=	VN_out_sigd(311);
CN_in_sigd(2409)	<=	VN_out_sigd(311);
CN_in_sigd(2641)	<=	VN_out_sigd(311);
CN_in_sigd(4193)	<=	VN_out_sigd(311);
CN_in_sigd(521)	<=	VN_out_sigd(312);
CN_in_sigd(2417)	<=	VN_out_sigd(312);
CN_in_sigd(2649)	<=	VN_out_sigd(312);
CN_in_sigd(4201)	<=	VN_out_sigd(312);
CN_in_sigd(529)	<=	VN_out_sigd(313);
CN_in_sigd(2425)	<=	VN_out_sigd(313);
CN_in_sigd(2657)	<=	VN_out_sigd(313);
CN_in_sigd(4209)	<=	VN_out_sigd(313);
CN_in_sigd(537)	<=	VN_out_sigd(314);
CN_in_sigd(2433)	<=	VN_out_sigd(314);
CN_in_sigd(2665)	<=	VN_out_sigd(314);
CN_in_sigd(4217)	<=	VN_out_sigd(314);
CN_in_sigd(545)	<=	VN_out_sigd(315);
CN_in_sigd(2441)	<=	VN_out_sigd(315);
CN_in_sigd(2673)	<=	VN_out_sigd(315);
CN_in_sigd(4225)	<=	VN_out_sigd(315);
CN_in_sigd(553)	<=	VN_out_sigd(316);
CN_in_sigd(2449)	<=	VN_out_sigd(316);
CN_in_sigd(2681)	<=	VN_out_sigd(316);
CN_in_sigd(4233)	<=	VN_out_sigd(316);
CN_in_sigd(561)	<=	VN_out_sigd(317);
CN_in_sigd(2457)	<=	VN_out_sigd(317);
CN_in_sigd(2689)	<=	VN_out_sigd(317);
CN_in_sigd(4241)	<=	VN_out_sigd(317);
CN_in_sigd(569)	<=	VN_out_sigd(318);
CN_in_sigd(2465)	<=	VN_out_sigd(318);
CN_in_sigd(2697)	<=	VN_out_sigd(318);
CN_in_sigd(4249)	<=	VN_out_sigd(318);
CN_in_sigd(577)	<=	VN_out_sigd(319);
CN_in_sigd(2473)	<=	VN_out_sigd(319);
CN_in_sigd(2705)	<=	VN_out_sigd(319);
CN_in_sigd(4257)	<=	VN_out_sigd(319);
CN_in_sigd(585)	<=	VN_out_sigd(320);
CN_in_sigd(2481)	<=	VN_out_sigd(320);
CN_in_sigd(2713)	<=	VN_out_sigd(320);
CN_in_sigd(4265)	<=	VN_out_sigd(320);
CN_in_sigd(593)	<=	VN_out_sigd(321);
CN_in_sigd(2489)	<=	VN_out_sigd(321);
CN_in_sigd(2721)	<=	VN_out_sigd(321);
CN_in_sigd(4273)	<=	VN_out_sigd(321);
CN_in_sigd(601)	<=	VN_out_sigd(322);
CN_in_sigd(2497)	<=	VN_out_sigd(322);
CN_in_sigd(2729)	<=	VN_out_sigd(322);
CN_in_sigd(4281)	<=	VN_out_sigd(322);
CN_in_sigd(609)	<=	VN_out_sigd(323);
CN_in_sigd(2505)	<=	VN_out_sigd(323);
CN_in_sigd(2737)	<=	VN_out_sigd(323);
CN_in_sigd(4289)	<=	VN_out_sigd(323);
CN_in_sigd(634)	<=	VN_out_sigd(324);
CN_in_sigd(1570)	<=	VN_out_sigd(324);
CN_in_sigd(3730)	<=	VN_out_sigd(324);
CN_in_sigd(4898)	<=	VN_out_sigd(324);
CN_in_sigd(642)	<=	VN_out_sigd(325);
CN_in_sigd(1578)	<=	VN_out_sigd(325);
CN_in_sigd(3738)	<=	VN_out_sigd(325);
CN_in_sigd(4906)	<=	VN_out_sigd(325);
CN_in_sigd(650)	<=	VN_out_sigd(326);
CN_in_sigd(1586)	<=	VN_out_sigd(326);
CN_in_sigd(3746)	<=	VN_out_sigd(326);
CN_in_sigd(4914)	<=	VN_out_sigd(326);
CN_in_sigd(658)	<=	VN_out_sigd(327);
CN_in_sigd(1594)	<=	VN_out_sigd(327);
CN_in_sigd(3754)	<=	VN_out_sigd(327);
CN_in_sigd(4922)	<=	VN_out_sigd(327);
CN_in_sigd(666)	<=	VN_out_sigd(328);
CN_in_sigd(1602)	<=	VN_out_sigd(328);
CN_in_sigd(3762)	<=	VN_out_sigd(328);
CN_in_sigd(4930)	<=	VN_out_sigd(328);
CN_in_sigd(674)	<=	VN_out_sigd(329);
CN_in_sigd(1610)	<=	VN_out_sigd(329);
CN_in_sigd(3770)	<=	VN_out_sigd(329);
CN_in_sigd(4938)	<=	VN_out_sigd(329);
CN_in_sigd(682)	<=	VN_out_sigd(330);
CN_in_sigd(1618)	<=	VN_out_sigd(330);
CN_in_sigd(3778)	<=	VN_out_sigd(330);
CN_in_sigd(4946)	<=	VN_out_sigd(330);
CN_in_sigd(690)	<=	VN_out_sigd(331);
CN_in_sigd(1626)	<=	VN_out_sigd(331);
CN_in_sigd(3786)	<=	VN_out_sigd(331);
CN_in_sigd(4954)	<=	VN_out_sigd(331);
CN_in_sigd(698)	<=	VN_out_sigd(332);
CN_in_sigd(1634)	<=	VN_out_sigd(332);
CN_in_sigd(3794)	<=	VN_out_sigd(332);
CN_in_sigd(4962)	<=	VN_out_sigd(332);
CN_in_sigd(706)	<=	VN_out_sigd(333);
CN_in_sigd(1642)	<=	VN_out_sigd(333);
CN_in_sigd(3802)	<=	VN_out_sigd(333);
CN_in_sigd(4970)	<=	VN_out_sigd(333);
CN_in_sigd(714)	<=	VN_out_sigd(334);
CN_in_sigd(1650)	<=	VN_out_sigd(334);
CN_in_sigd(3810)	<=	VN_out_sigd(334);
CN_in_sigd(4978)	<=	VN_out_sigd(334);
CN_in_sigd(722)	<=	VN_out_sigd(335);
CN_in_sigd(1658)	<=	VN_out_sigd(335);
CN_in_sigd(3818)	<=	VN_out_sigd(335);
CN_in_sigd(4986)	<=	VN_out_sigd(335);
CN_in_sigd(730)	<=	VN_out_sigd(336);
CN_in_sigd(1666)	<=	VN_out_sigd(336);
CN_in_sigd(3826)	<=	VN_out_sigd(336);
CN_in_sigd(4994)	<=	VN_out_sigd(336);
CN_in_sigd(738)	<=	VN_out_sigd(337);
CN_in_sigd(1674)	<=	VN_out_sigd(337);
CN_in_sigd(3834)	<=	VN_out_sigd(337);
CN_in_sigd(5002)	<=	VN_out_sigd(337);
CN_in_sigd(746)	<=	VN_out_sigd(338);
CN_in_sigd(1682)	<=	VN_out_sigd(338);
CN_in_sigd(3842)	<=	VN_out_sigd(338);
CN_in_sigd(5010)	<=	VN_out_sigd(338);
CN_in_sigd(754)	<=	VN_out_sigd(339);
CN_in_sigd(1690)	<=	VN_out_sigd(339);
CN_in_sigd(3850)	<=	VN_out_sigd(339);
CN_in_sigd(5018)	<=	VN_out_sigd(339);
CN_in_sigd(762)	<=	VN_out_sigd(340);
CN_in_sigd(1698)	<=	VN_out_sigd(340);
CN_in_sigd(3858)	<=	VN_out_sigd(340);
CN_in_sigd(5026)	<=	VN_out_sigd(340);
CN_in_sigd(770)	<=	VN_out_sigd(341);
CN_in_sigd(1706)	<=	VN_out_sigd(341);
CN_in_sigd(3866)	<=	VN_out_sigd(341);
CN_in_sigd(5034)	<=	VN_out_sigd(341);
CN_in_sigd(778)	<=	VN_out_sigd(342);
CN_in_sigd(1714)	<=	VN_out_sigd(342);
CN_in_sigd(3874)	<=	VN_out_sigd(342);
CN_in_sigd(5042)	<=	VN_out_sigd(342);
CN_in_sigd(786)	<=	VN_out_sigd(343);
CN_in_sigd(1722)	<=	VN_out_sigd(343);
CN_in_sigd(3882)	<=	VN_out_sigd(343);
CN_in_sigd(5050)	<=	VN_out_sigd(343);
CN_in_sigd(794)	<=	VN_out_sigd(344);
CN_in_sigd(1298)	<=	VN_out_sigd(344);
CN_in_sigd(3458)	<=	VN_out_sigd(344);
CN_in_sigd(5058)	<=	VN_out_sigd(344);
CN_in_sigd(802)	<=	VN_out_sigd(345);
CN_in_sigd(1306)	<=	VN_out_sigd(345);
CN_in_sigd(3466)	<=	VN_out_sigd(345);
CN_in_sigd(5066)	<=	VN_out_sigd(345);
CN_in_sigd(810)	<=	VN_out_sigd(346);
CN_in_sigd(1314)	<=	VN_out_sigd(346);
CN_in_sigd(3474)	<=	VN_out_sigd(346);
CN_in_sigd(5074)	<=	VN_out_sigd(346);
CN_in_sigd(818)	<=	VN_out_sigd(347);
CN_in_sigd(1322)	<=	VN_out_sigd(347);
CN_in_sigd(3482)	<=	VN_out_sigd(347);
CN_in_sigd(5082)	<=	VN_out_sigd(347);
CN_in_sigd(826)	<=	VN_out_sigd(348);
CN_in_sigd(1330)	<=	VN_out_sigd(348);
CN_in_sigd(3490)	<=	VN_out_sigd(348);
CN_in_sigd(5090)	<=	VN_out_sigd(348);
CN_in_sigd(834)	<=	VN_out_sigd(349);
CN_in_sigd(1338)	<=	VN_out_sigd(349);
CN_in_sigd(3498)	<=	VN_out_sigd(349);
CN_in_sigd(5098)	<=	VN_out_sigd(349);
CN_in_sigd(842)	<=	VN_out_sigd(350);
CN_in_sigd(1346)	<=	VN_out_sigd(350);
CN_in_sigd(3506)	<=	VN_out_sigd(350);
CN_in_sigd(5106)	<=	VN_out_sigd(350);
CN_in_sigd(850)	<=	VN_out_sigd(351);
CN_in_sigd(1354)	<=	VN_out_sigd(351);
CN_in_sigd(3514)	<=	VN_out_sigd(351);
CN_in_sigd(5114)	<=	VN_out_sigd(351);
CN_in_sigd(858)	<=	VN_out_sigd(352);
CN_in_sigd(1362)	<=	VN_out_sigd(352);
CN_in_sigd(3522)	<=	VN_out_sigd(352);
CN_in_sigd(5122)	<=	VN_out_sigd(352);
CN_in_sigd(434)	<=	VN_out_sigd(353);
CN_in_sigd(1370)	<=	VN_out_sigd(353);
CN_in_sigd(3530)	<=	VN_out_sigd(353);
CN_in_sigd(5130)	<=	VN_out_sigd(353);
CN_in_sigd(442)	<=	VN_out_sigd(354);
CN_in_sigd(1378)	<=	VN_out_sigd(354);
CN_in_sigd(3538)	<=	VN_out_sigd(354);
CN_in_sigd(5138)	<=	VN_out_sigd(354);
CN_in_sigd(450)	<=	VN_out_sigd(355);
CN_in_sigd(1386)	<=	VN_out_sigd(355);
CN_in_sigd(3546)	<=	VN_out_sigd(355);
CN_in_sigd(5146)	<=	VN_out_sigd(355);
CN_in_sigd(458)	<=	VN_out_sigd(356);
CN_in_sigd(1394)	<=	VN_out_sigd(356);
CN_in_sigd(3554)	<=	VN_out_sigd(356);
CN_in_sigd(5154)	<=	VN_out_sigd(356);
CN_in_sigd(466)	<=	VN_out_sigd(357);
CN_in_sigd(1402)	<=	VN_out_sigd(357);
CN_in_sigd(3562)	<=	VN_out_sigd(357);
CN_in_sigd(5162)	<=	VN_out_sigd(357);
CN_in_sigd(474)	<=	VN_out_sigd(358);
CN_in_sigd(1410)	<=	VN_out_sigd(358);
CN_in_sigd(3570)	<=	VN_out_sigd(358);
CN_in_sigd(5170)	<=	VN_out_sigd(358);
CN_in_sigd(482)	<=	VN_out_sigd(359);
CN_in_sigd(1418)	<=	VN_out_sigd(359);
CN_in_sigd(3578)	<=	VN_out_sigd(359);
CN_in_sigd(5178)	<=	VN_out_sigd(359);
CN_in_sigd(490)	<=	VN_out_sigd(360);
CN_in_sigd(1426)	<=	VN_out_sigd(360);
CN_in_sigd(3586)	<=	VN_out_sigd(360);
CN_in_sigd(4754)	<=	VN_out_sigd(360);
CN_in_sigd(498)	<=	VN_out_sigd(361);
CN_in_sigd(1434)	<=	VN_out_sigd(361);
CN_in_sigd(3594)	<=	VN_out_sigd(361);
CN_in_sigd(4762)	<=	VN_out_sigd(361);
CN_in_sigd(506)	<=	VN_out_sigd(362);
CN_in_sigd(1442)	<=	VN_out_sigd(362);
CN_in_sigd(3602)	<=	VN_out_sigd(362);
CN_in_sigd(4770)	<=	VN_out_sigd(362);
CN_in_sigd(514)	<=	VN_out_sigd(363);
CN_in_sigd(1450)	<=	VN_out_sigd(363);
CN_in_sigd(3610)	<=	VN_out_sigd(363);
CN_in_sigd(4778)	<=	VN_out_sigd(363);
CN_in_sigd(522)	<=	VN_out_sigd(364);
CN_in_sigd(1458)	<=	VN_out_sigd(364);
CN_in_sigd(3618)	<=	VN_out_sigd(364);
CN_in_sigd(4786)	<=	VN_out_sigd(364);
CN_in_sigd(530)	<=	VN_out_sigd(365);
CN_in_sigd(1466)	<=	VN_out_sigd(365);
CN_in_sigd(3626)	<=	VN_out_sigd(365);
CN_in_sigd(4794)	<=	VN_out_sigd(365);
CN_in_sigd(538)	<=	VN_out_sigd(366);
CN_in_sigd(1474)	<=	VN_out_sigd(366);
CN_in_sigd(3634)	<=	VN_out_sigd(366);
CN_in_sigd(4802)	<=	VN_out_sigd(366);
CN_in_sigd(546)	<=	VN_out_sigd(367);
CN_in_sigd(1482)	<=	VN_out_sigd(367);
CN_in_sigd(3642)	<=	VN_out_sigd(367);
CN_in_sigd(4810)	<=	VN_out_sigd(367);
CN_in_sigd(554)	<=	VN_out_sigd(368);
CN_in_sigd(1490)	<=	VN_out_sigd(368);
CN_in_sigd(3650)	<=	VN_out_sigd(368);
CN_in_sigd(4818)	<=	VN_out_sigd(368);
CN_in_sigd(562)	<=	VN_out_sigd(369);
CN_in_sigd(1498)	<=	VN_out_sigd(369);
CN_in_sigd(3658)	<=	VN_out_sigd(369);
CN_in_sigd(4826)	<=	VN_out_sigd(369);
CN_in_sigd(570)	<=	VN_out_sigd(370);
CN_in_sigd(1506)	<=	VN_out_sigd(370);
CN_in_sigd(3666)	<=	VN_out_sigd(370);
CN_in_sigd(4834)	<=	VN_out_sigd(370);
CN_in_sigd(578)	<=	VN_out_sigd(371);
CN_in_sigd(1514)	<=	VN_out_sigd(371);
CN_in_sigd(3674)	<=	VN_out_sigd(371);
CN_in_sigd(4842)	<=	VN_out_sigd(371);
CN_in_sigd(586)	<=	VN_out_sigd(372);
CN_in_sigd(1522)	<=	VN_out_sigd(372);
CN_in_sigd(3682)	<=	VN_out_sigd(372);
CN_in_sigd(4850)	<=	VN_out_sigd(372);
CN_in_sigd(594)	<=	VN_out_sigd(373);
CN_in_sigd(1530)	<=	VN_out_sigd(373);
CN_in_sigd(3690)	<=	VN_out_sigd(373);
CN_in_sigd(4858)	<=	VN_out_sigd(373);
CN_in_sigd(602)	<=	VN_out_sigd(374);
CN_in_sigd(1538)	<=	VN_out_sigd(374);
CN_in_sigd(3698)	<=	VN_out_sigd(374);
CN_in_sigd(4866)	<=	VN_out_sigd(374);
CN_in_sigd(610)	<=	VN_out_sigd(375);
CN_in_sigd(1546)	<=	VN_out_sigd(375);
CN_in_sigd(3706)	<=	VN_out_sigd(375);
CN_in_sigd(4874)	<=	VN_out_sigd(375);
CN_in_sigd(618)	<=	VN_out_sigd(376);
CN_in_sigd(1554)	<=	VN_out_sigd(376);
CN_in_sigd(3714)	<=	VN_out_sigd(376);
CN_in_sigd(4882)	<=	VN_out_sigd(376);
CN_in_sigd(626)	<=	VN_out_sigd(377);
CN_in_sigd(1562)	<=	VN_out_sigd(377);
CN_in_sigd(3722)	<=	VN_out_sigd(377);
CN_in_sigd(4890)	<=	VN_out_sigd(377);
CN_in_sigd(1210)	<=	VN_out_sigd(378);
CN_in_sigd(2074)	<=	VN_out_sigd(378);
CN_in_sigd(3226)	<=	VN_out_sigd(378);
CN_in_sigd(4714)	<=	VN_out_sigd(378);
CN_in_sigd(1218)	<=	VN_out_sigd(379);
CN_in_sigd(2082)	<=	VN_out_sigd(379);
CN_in_sigd(3234)	<=	VN_out_sigd(379);
CN_in_sigd(4722)	<=	VN_out_sigd(379);
CN_in_sigd(1226)	<=	VN_out_sigd(380);
CN_in_sigd(2090)	<=	VN_out_sigd(380);
CN_in_sigd(3242)	<=	VN_out_sigd(380);
CN_in_sigd(4730)	<=	VN_out_sigd(380);
CN_in_sigd(1234)	<=	VN_out_sigd(381);
CN_in_sigd(2098)	<=	VN_out_sigd(381);
CN_in_sigd(3250)	<=	VN_out_sigd(381);
CN_in_sigd(4738)	<=	VN_out_sigd(381);
CN_in_sigd(1242)	<=	VN_out_sigd(382);
CN_in_sigd(2106)	<=	VN_out_sigd(382);
CN_in_sigd(3258)	<=	VN_out_sigd(382);
CN_in_sigd(4746)	<=	VN_out_sigd(382);
CN_in_sigd(1250)	<=	VN_out_sigd(383);
CN_in_sigd(2114)	<=	VN_out_sigd(383);
CN_in_sigd(3266)	<=	VN_out_sigd(383);
CN_in_sigd(4322)	<=	VN_out_sigd(383);
CN_in_sigd(1258)	<=	VN_out_sigd(384);
CN_in_sigd(2122)	<=	VN_out_sigd(384);
CN_in_sigd(3274)	<=	VN_out_sigd(384);
CN_in_sigd(4330)	<=	VN_out_sigd(384);
CN_in_sigd(1266)	<=	VN_out_sigd(385);
CN_in_sigd(2130)	<=	VN_out_sigd(385);
CN_in_sigd(3282)	<=	VN_out_sigd(385);
CN_in_sigd(4338)	<=	VN_out_sigd(385);
CN_in_sigd(1274)	<=	VN_out_sigd(386);
CN_in_sigd(2138)	<=	VN_out_sigd(386);
CN_in_sigd(3290)	<=	VN_out_sigd(386);
CN_in_sigd(4346)	<=	VN_out_sigd(386);
CN_in_sigd(1282)	<=	VN_out_sigd(387);
CN_in_sigd(2146)	<=	VN_out_sigd(387);
CN_in_sigd(3298)	<=	VN_out_sigd(387);
CN_in_sigd(4354)	<=	VN_out_sigd(387);
CN_in_sigd(1290)	<=	VN_out_sigd(388);
CN_in_sigd(2154)	<=	VN_out_sigd(388);
CN_in_sigd(3306)	<=	VN_out_sigd(388);
CN_in_sigd(4362)	<=	VN_out_sigd(388);
CN_in_sigd(866)	<=	VN_out_sigd(389);
CN_in_sigd(1730)	<=	VN_out_sigd(389);
CN_in_sigd(3314)	<=	VN_out_sigd(389);
CN_in_sigd(4370)	<=	VN_out_sigd(389);
CN_in_sigd(874)	<=	VN_out_sigd(390);
CN_in_sigd(1738)	<=	VN_out_sigd(390);
CN_in_sigd(3322)	<=	VN_out_sigd(390);
CN_in_sigd(4378)	<=	VN_out_sigd(390);
CN_in_sigd(882)	<=	VN_out_sigd(391);
CN_in_sigd(1746)	<=	VN_out_sigd(391);
CN_in_sigd(3330)	<=	VN_out_sigd(391);
CN_in_sigd(4386)	<=	VN_out_sigd(391);
CN_in_sigd(890)	<=	VN_out_sigd(392);
CN_in_sigd(1754)	<=	VN_out_sigd(392);
CN_in_sigd(3338)	<=	VN_out_sigd(392);
CN_in_sigd(4394)	<=	VN_out_sigd(392);
CN_in_sigd(898)	<=	VN_out_sigd(393);
CN_in_sigd(1762)	<=	VN_out_sigd(393);
CN_in_sigd(3346)	<=	VN_out_sigd(393);
CN_in_sigd(4402)	<=	VN_out_sigd(393);
CN_in_sigd(906)	<=	VN_out_sigd(394);
CN_in_sigd(1770)	<=	VN_out_sigd(394);
CN_in_sigd(3354)	<=	VN_out_sigd(394);
CN_in_sigd(4410)	<=	VN_out_sigd(394);
CN_in_sigd(914)	<=	VN_out_sigd(395);
CN_in_sigd(1778)	<=	VN_out_sigd(395);
CN_in_sigd(3362)	<=	VN_out_sigd(395);
CN_in_sigd(4418)	<=	VN_out_sigd(395);
CN_in_sigd(922)	<=	VN_out_sigd(396);
CN_in_sigd(1786)	<=	VN_out_sigd(396);
CN_in_sigd(3370)	<=	VN_out_sigd(396);
CN_in_sigd(4426)	<=	VN_out_sigd(396);
CN_in_sigd(930)	<=	VN_out_sigd(397);
CN_in_sigd(1794)	<=	VN_out_sigd(397);
CN_in_sigd(3378)	<=	VN_out_sigd(397);
CN_in_sigd(4434)	<=	VN_out_sigd(397);
CN_in_sigd(938)	<=	VN_out_sigd(398);
CN_in_sigd(1802)	<=	VN_out_sigd(398);
CN_in_sigd(3386)	<=	VN_out_sigd(398);
CN_in_sigd(4442)	<=	VN_out_sigd(398);
CN_in_sigd(946)	<=	VN_out_sigd(399);
CN_in_sigd(1810)	<=	VN_out_sigd(399);
CN_in_sigd(3394)	<=	VN_out_sigd(399);
CN_in_sigd(4450)	<=	VN_out_sigd(399);
CN_in_sigd(954)	<=	VN_out_sigd(400);
CN_in_sigd(1818)	<=	VN_out_sigd(400);
CN_in_sigd(3402)	<=	VN_out_sigd(400);
CN_in_sigd(4458)	<=	VN_out_sigd(400);
CN_in_sigd(962)	<=	VN_out_sigd(401);
CN_in_sigd(1826)	<=	VN_out_sigd(401);
CN_in_sigd(3410)	<=	VN_out_sigd(401);
CN_in_sigd(4466)	<=	VN_out_sigd(401);
CN_in_sigd(970)	<=	VN_out_sigd(402);
CN_in_sigd(1834)	<=	VN_out_sigd(402);
CN_in_sigd(3418)	<=	VN_out_sigd(402);
CN_in_sigd(4474)	<=	VN_out_sigd(402);
CN_in_sigd(978)	<=	VN_out_sigd(403);
CN_in_sigd(1842)	<=	VN_out_sigd(403);
CN_in_sigd(3426)	<=	VN_out_sigd(403);
CN_in_sigd(4482)	<=	VN_out_sigd(403);
CN_in_sigd(986)	<=	VN_out_sigd(404);
CN_in_sigd(1850)	<=	VN_out_sigd(404);
CN_in_sigd(3434)	<=	VN_out_sigd(404);
CN_in_sigd(4490)	<=	VN_out_sigd(404);
CN_in_sigd(994)	<=	VN_out_sigd(405);
CN_in_sigd(1858)	<=	VN_out_sigd(405);
CN_in_sigd(3442)	<=	VN_out_sigd(405);
CN_in_sigd(4498)	<=	VN_out_sigd(405);
CN_in_sigd(1002)	<=	VN_out_sigd(406);
CN_in_sigd(1866)	<=	VN_out_sigd(406);
CN_in_sigd(3450)	<=	VN_out_sigd(406);
CN_in_sigd(4506)	<=	VN_out_sigd(406);
CN_in_sigd(1010)	<=	VN_out_sigd(407);
CN_in_sigd(1874)	<=	VN_out_sigd(407);
CN_in_sigd(3026)	<=	VN_out_sigd(407);
CN_in_sigd(4514)	<=	VN_out_sigd(407);
CN_in_sigd(1018)	<=	VN_out_sigd(408);
CN_in_sigd(1882)	<=	VN_out_sigd(408);
CN_in_sigd(3034)	<=	VN_out_sigd(408);
CN_in_sigd(4522)	<=	VN_out_sigd(408);
CN_in_sigd(1026)	<=	VN_out_sigd(409);
CN_in_sigd(1890)	<=	VN_out_sigd(409);
CN_in_sigd(3042)	<=	VN_out_sigd(409);
CN_in_sigd(4530)	<=	VN_out_sigd(409);
CN_in_sigd(1034)	<=	VN_out_sigd(410);
CN_in_sigd(1898)	<=	VN_out_sigd(410);
CN_in_sigd(3050)	<=	VN_out_sigd(410);
CN_in_sigd(4538)	<=	VN_out_sigd(410);
CN_in_sigd(1042)	<=	VN_out_sigd(411);
CN_in_sigd(1906)	<=	VN_out_sigd(411);
CN_in_sigd(3058)	<=	VN_out_sigd(411);
CN_in_sigd(4546)	<=	VN_out_sigd(411);
CN_in_sigd(1050)	<=	VN_out_sigd(412);
CN_in_sigd(1914)	<=	VN_out_sigd(412);
CN_in_sigd(3066)	<=	VN_out_sigd(412);
CN_in_sigd(4554)	<=	VN_out_sigd(412);
CN_in_sigd(1058)	<=	VN_out_sigd(413);
CN_in_sigd(1922)	<=	VN_out_sigd(413);
CN_in_sigd(3074)	<=	VN_out_sigd(413);
CN_in_sigd(4562)	<=	VN_out_sigd(413);
CN_in_sigd(1066)	<=	VN_out_sigd(414);
CN_in_sigd(1930)	<=	VN_out_sigd(414);
CN_in_sigd(3082)	<=	VN_out_sigd(414);
CN_in_sigd(4570)	<=	VN_out_sigd(414);
CN_in_sigd(1074)	<=	VN_out_sigd(415);
CN_in_sigd(1938)	<=	VN_out_sigd(415);
CN_in_sigd(3090)	<=	VN_out_sigd(415);
CN_in_sigd(4578)	<=	VN_out_sigd(415);
CN_in_sigd(1082)	<=	VN_out_sigd(416);
CN_in_sigd(1946)	<=	VN_out_sigd(416);
CN_in_sigd(3098)	<=	VN_out_sigd(416);
CN_in_sigd(4586)	<=	VN_out_sigd(416);
CN_in_sigd(1090)	<=	VN_out_sigd(417);
CN_in_sigd(1954)	<=	VN_out_sigd(417);
CN_in_sigd(3106)	<=	VN_out_sigd(417);
CN_in_sigd(4594)	<=	VN_out_sigd(417);
CN_in_sigd(1098)	<=	VN_out_sigd(418);
CN_in_sigd(1962)	<=	VN_out_sigd(418);
CN_in_sigd(3114)	<=	VN_out_sigd(418);
CN_in_sigd(4602)	<=	VN_out_sigd(418);
CN_in_sigd(1106)	<=	VN_out_sigd(419);
CN_in_sigd(1970)	<=	VN_out_sigd(419);
CN_in_sigd(3122)	<=	VN_out_sigd(419);
CN_in_sigd(4610)	<=	VN_out_sigd(419);
CN_in_sigd(1114)	<=	VN_out_sigd(420);
CN_in_sigd(1978)	<=	VN_out_sigd(420);
CN_in_sigd(3130)	<=	VN_out_sigd(420);
CN_in_sigd(4618)	<=	VN_out_sigd(420);
CN_in_sigd(1122)	<=	VN_out_sigd(421);
CN_in_sigd(1986)	<=	VN_out_sigd(421);
CN_in_sigd(3138)	<=	VN_out_sigd(421);
CN_in_sigd(4626)	<=	VN_out_sigd(421);
CN_in_sigd(1130)	<=	VN_out_sigd(422);
CN_in_sigd(1994)	<=	VN_out_sigd(422);
CN_in_sigd(3146)	<=	VN_out_sigd(422);
CN_in_sigd(4634)	<=	VN_out_sigd(422);
CN_in_sigd(1138)	<=	VN_out_sigd(423);
CN_in_sigd(2002)	<=	VN_out_sigd(423);
CN_in_sigd(3154)	<=	VN_out_sigd(423);
CN_in_sigd(4642)	<=	VN_out_sigd(423);
CN_in_sigd(1146)	<=	VN_out_sigd(424);
CN_in_sigd(2010)	<=	VN_out_sigd(424);
CN_in_sigd(3162)	<=	VN_out_sigd(424);
CN_in_sigd(4650)	<=	VN_out_sigd(424);
CN_in_sigd(1154)	<=	VN_out_sigd(425);
CN_in_sigd(2018)	<=	VN_out_sigd(425);
CN_in_sigd(3170)	<=	VN_out_sigd(425);
CN_in_sigd(4658)	<=	VN_out_sigd(425);
CN_in_sigd(1162)	<=	VN_out_sigd(426);
CN_in_sigd(2026)	<=	VN_out_sigd(426);
CN_in_sigd(3178)	<=	VN_out_sigd(426);
CN_in_sigd(4666)	<=	VN_out_sigd(426);
CN_in_sigd(1170)	<=	VN_out_sigd(427);
CN_in_sigd(2034)	<=	VN_out_sigd(427);
CN_in_sigd(3186)	<=	VN_out_sigd(427);
CN_in_sigd(4674)	<=	VN_out_sigd(427);
CN_in_sigd(1178)	<=	VN_out_sigd(428);
CN_in_sigd(2042)	<=	VN_out_sigd(428);
CN_in_sigd(3194)	<=	VN_out_sigd(428);
CN_in_sigd(4682)	<=	VN_out_sigd(428);
CN_in_sigd(1186)	<=	VN_out_sigd(429);
CN_in_sigd(2050)	<=	VN_out_sigd(429);
CN_in_sigd(3202)	<=	VN_out_sigd(429);
CN_in_sigd(4690)	<=	VN_out_sigd(429);
CN_in_sigd(1194)	<=	VN_out_sigd(430);
CN_in_sigd(2058)	<=	VN_out_sigd(430);
CN_in_sigd(3210)	<=	VN_out_sigd(430);
CN_in_sigd(4698)	<=	VN_out_sigd(430);
CN_in_sigd(1202)	<=	VN_out_sigd(431);
CN_in_sigd(2066)	<=	VN_out_sigd(431);
CN_in_sigd(3218)	<=	VN_out_sigd(431);
CN_in_sigd(4706)	<=	VN_out_sigd(431);
CN_in_sigd(170)	<=	VN_out_sigd(432);
CN_in_sigd(2514)	<=	VN_out_sigd(432);
CN_in_sigd(2778)	<=	VN_out_sigd(432);
CN_in_sigd(4114)	<=	VN_out_sigd(432);
CN_in_sigd(178)	<=	VN_out_sigd(433);
CN_in_sigd(2522)	<=	VN_out_sigd(433);
CN_in_sigd(2786)	<=	VN_out_sigd(433);
CN_in_sigd(4122)	<=	VN_out_sigd(433);
CN_in_sigd(186)	<=	VN_out_sigd(434);
CN_in_sigd(2530)	<=	VN_out_sigd(434);
CN_in_sigd(2794)	<=	VN_out_sigd(434);
CN_in_sigd(4130)	<=	VN_out_sigd(434);
CN_in_sigd(194)	<=	VN_out_sigd(435);
CN_in_sigd(2538)	<=	VN_out_sigd(435);
CN_in_sigd(2802)	<=	VN_out_sigd(435);
CN_in_sigd(4138)	<=	VN_out_sigd(435);
CN_in_sigd(202)	<=	VN_out_sigd(436);
CN_in_sigd(2546)	<=	VN_out_sigd(436);
CN_in_sigd(2810)	<=	VN_out_sigd(436);
CN_in_sigd(4146)	<=	VN_out_sigd(436);
CN_in_sigd(210)	<=	VN_out_sigd(437);
CN_in_sigd(2554)	<=	VN_out_sigd(437);
CN_in_sigd(2818)	<=	VN_out_sigd(437);
CN_in_sigd(4154)	<=	VN_out_sigd(437);
CN_in_sigd(218)	<=	VN_out_sigd(438);
CN_in_sigd(2562)	<=	VN_out_sigd(438);
CN_in_sigd(2826)	<=	VN_out_sigd(438);
CN_in_sigd(4162)	<=	VN_out_sigd(438);
CN_in_sigd(226)	<=	VN_out_sigd(439);
CN_in_sigd(2570)	<=	VN_out_sigd(439);
CN_in_sigd(2834)	<=	VN_out_sigd(439);
CN_in_sigd(4170)	<=	VN_out_sigd(439);
CN_in_sigd(234)	<=	VN_out_sigd(440);
CN_in_sigd(2578)	<=	VN_out_sigd(440);
CN_in_sigd(2842)	<=	VN_out_sigd(440);
CN_in_sigd(4178)	<=	VN_out_sigd(440);
CN_in_sigd(242)	<=	VN_out_sigd(441);
CN_in_sigd(2586)	<=	VN_out_sigd(441);
CN_in_sigd(2850)	<=	VN_out_sigd(441);
CN_in_sigd(4186)	<=	VN_out_sigd(441);
CN_in_sigd(250)	<=	VN_out_sigd(442);
CN_in_sigd(2162)	<=	VN_out_sigd(442);
CN_in_sigd(2858)	<=	VN_out_sigd(442);
CN_in_sigd(4194)	<=	VN_out_sigd(442);
CN_in_sigd(258)	<=	VN_out_sigd(443);
CN_in_sigd(2170)	<=	VN_out_sigd(443);
CN_in_sigd(2866)	<=	VN_out_sigd(443);
CN_in_sigd(4202)	<=	VN_out_sigd(443);
CN_in_sigd(266)	<=	VN_out_sigd(444);
CN_in_sigd(2178)	<=	VN_out_sigd(444);
CN_in_sigd(2874)	<=	VN_out_sigd(444);
CN_in_sigd(4210)	<=	VN_out_sigd(444);
CN_in_sigd(274)	<=	VN_out_sigd(445);
CN_in_sigd(2186)	<=	VN_out_sigd(445);
CN_in_sigd(2882)	<=	VN_out_sigd(445);
CN_in_sigd(4218)	<=	VN_out_sigd(445);
CN_in_sigd(282)	<=	VN_out_sigd(446);
CN_in_sigd(2194)	<=	VN_out_sigd(446);
CN_in_sigd(2890)	<=	VN_out_sigd(446);
CN_in_sigd(4226)	<=	VN_out_sigd(446);
CN_in_sigd(290)	<=	VN_out_sigd(447);
CN_in_sigd(2202)	<=	VN_out_sigd(447);
CN_in_sigd(2898)	<=	VN_out_sigd(447);
CN_in_sigd(4234)	<=	VN_out_sigd(447);
CN_in_sigd(298)	<=	VN_out_sigd(448);
CN_in_sigd(2210)	<=	VN_out_sigd(448);
CN_in_sigd(2906)	<=	VN_out_sigd(448);
CN_in_sigd(4242)	<=	VN_out_sigd(448);
CN_in_sigd(306)	<=	VN_out_sigd(449);
CN_in_sigd(2218)	<=	VN_out_sigd(449);
CN_in_sigd(2914)	<=	VN_out_sigd(449);
CN_in_sigd(4250)	<=	VN_out_sigd(449);
CN_in_sigd(314)	<=	VN_out_sigd(450);
CN_in_sigd(2226)	<=	VN_out_sigd(450);
CN_in_sigd(2922)	<=	VN_out_sigd(450);
CN_in_sigd(4258)	<=	VN_out_sigd(450);
CN_in_sigd(322)	<=	VN_out_sigd(451);
CN_in_sigd(2234)	<=	VN_out_sigd(451);
CN_in_sigd(2930)	<=	VN_out_sigd(451);
CN_in_sigd(4266)	<=	VN_out_sigd(451);
CN_in_sigd(330)	<=	VN_out_sigd(452);
CN_in_sigd(2242)	<=	VN_out_sigd(452);
CN_in_sigd(2938)	<=	VN_out_sigd(452);
CN_in_sigd(4274)	<=	VN_out_sigd(452);
CN_in_sigd(338)	<=	VN_out_sigd(453);
CN_in_sigd(2250)	<=	VN_out_sigd(453);
CN_in_sigd(2946)	<=	VN_out_sigd(453);
CN_in_sigd(4282)	<=	VN_out_sigd(453);
CN_in_sigd(346)	<=	VN_out_sigd(454);
CN_in_sigd(2258)	<=	VN_out_sigd(454);
CN_in_sigd(2954)	<=	VN_out_sigd(454);
CN_in_sigd(4290)	<=	VN_out_sigd(454);
CN_in_sigd(354)	<=	VN_out_sigd(455);
CN_in_sigd(2266)	<=	VN_out_sigd(455);
CN_in_sigd(2962)	<=	VN_out_sigd(455);
CN_in_sigd(4298)	<=	VN_out_sigd(455);
CN_in_sigd(362)	<=	VN_out_sigd(456);
CN_in_sigd(2274)	<=	VN_out_sigd(456);
CN_in_sigd(2970)	<=	VN_out_sigd(456);
CN_in_sigd(4306)	<=	VN_out_sigd(456);
CN_in_sigd(370)	<=	VN_out_sigd(457);
CN_in_sigd(2282)	<=	VN_out_sigd(457);
CN_in_sigd(2978)	<=	VN_out_sigd(457);
CN_in_sigd(4314)	<=	VN_out_sigd(457);
CN_in_sigd(378)	<=	VN_out_sigd(458);
CN_in_sigd(2290)	<=	VN_out_sigd(458);
CN_in_sigd(2986)	<=	VN_out_sigd(458);
CN_in_sigd(3890)	<=	VN_out_sigd(458);
CN_in_sigd(386)	<=	VN_out_sigd(459);
CN_in_sigd(2298)	<=	VN_out_sigd(459);
CN_in_sigd(2994)	<=	VN_out_sigd(459);
CN_in_sigd(3898)	<=	VN_out_sigd(459);
CN_in_sigd(394)	<=	VN_out_sigd(460);
CN_in_sigd(2306)	<=	VN_out_sigd(460);
CN_in_sigd(3002)	<=	VN_out_sigd(460);
CN_in_sigd(3906)	<=	VN_out_sigd(460);
CN_in_sigd(402)	<=	VN_out_sigd(461);
CN_in_sigd(2314)	<=	VN_out_sigd(461);
CN_in_sigd(3010)	<=	VN_out_sigd(461);
CN_in_sigd(3914)	<=	VN_out_sigd(461);
CN_in_sigd(410)	<=	VN_out_sigd(462);
CN_in_sigd(2322)	<=	VN_out_sigd(462);
CN_in_sigd(3018)	<=	VN_out_sigd(462);
CN_in_sigd(3922)	<=	VN_out_sigd(462);
CN_in_sigd(418)	<=	VN_out_sigd(463);
CN_in_sigd(2330)	<=	VN_out_sigd(463);
CN_in_sigd(2594)	<=	VN_out_sigd(463);
CN_in_sigd(3930)	<=	VN_out_sigd(463);
CN_in_sigd(426)	<=	VN_out_sigd(464);
CN_in_sigd(2338)	<=	VN_out_sigd(464);
CN_in_sigd(2602)	<=	VN_out_sigd(464);
CN_in_sigd(3938)	<=	VN_out_sigd(464);
CN_in_sigd(2)	<=	VN_out_sigd(465);
CN_in_sigd(2346)	<=	VN_out_sigd(465);
CN_in_sigd(2610)	<=	VN_out_sigd(465);
CN_in_sigd(3946)	<=	VN_out_sigd(465);
CN_in_sigd(10)	<=	VN_out_sigd(466);
CN_in_sigd(2354)	<=	VN_out_sigd(466);
CN_in_sigd(2618)	<=	VN_out_sigd(466);
CN_in_sigd(3954)	<=	VN_out_sigd(466);
CN_in_sigd(18)	<=	VN_out_sigd(467);
CN_in_sigd(2362)	<=	VN_out_sigd(467);
CN_in_sigd(2626)	<=	VN_out_sigd(467);
CN_in_sigd(3962)	<=	VN_out_sigd(467);
CN_in_sigd(26)	<=	VN_out_sigd(468);
CN_in_sigd(2370)	<=	VN_out_sigd(468);
CN_in_sigd(2634)	<=	VN_out_sigd(468);
CN_in_sigd(3970)	<=	VN_out_sigd(468);
CN_in_sigd(34)	<=	VN_out_sigd(469);
CN_in_sigd(2378)	<=	VN_out_sigd(469);
CN_in_sigd(2642)	<=	VN_out_sigd(469);
CN_in_sigd(3978)	<=	VN_out_sigd(469);
CN_in_sigd(42)	<=	VN_out_sigd(470);
CN_in_sigd(2386)	<=	VN_out_sigd(470);
CN_in_sigd(2650)	<=	VN_out_sigd(470);
CN_in_sigd(3986)	<=	VN_out_sigd(470);
CN_in_sigd(50)	<=	VN_out_sigd(471);
CN_in_sigd(2394)	<=	VN_out_sigd(471);
CN_in_sigd(2658)	<=	VN_out_sigd(471);
CN_in_sigd(3994)	<=	VN_out_sigd(471);
CN_in_sigd(58)	<=	VN_out_sigd(472);
CN_in_sigd(2402)	<=	VN_out_sigd(472);
CN_in_sigd(2666)	<=	VN_out_sigd(472);
CN_in_sigd(4002)	<=	VN_out_sigd(472);
CN_in_sigd(66)	<=	VN_out_sigd(473);
CN_in_sigd(2410)	<=	VN_out_sigd(473);
CN_in_sigd(2674)	<=	VN_out_sigd(473);
CN_in_sigd(4010)	<=	VN_out_sigd(473);
CN_in_sigd(74)	<=	VN_out_sigd(474);
CN_in_sigd(2418)	<=	VN_out_sigd(474);
CN_in_sigd(2682)	<=	VN_out_sigd(474);
CN_in_sigd(4018)	<=	VN_out_sigd(474);
CN_in_sigd(82)	<=	VN_out_sigd(475);
CN_in_sigd(2426)	<=	VN_out_sigd(475);
CN_in_sigd(2690)	<=	VN_out_sigd(475);
CN_in_sigd(4026)	<=	VN_out_sigd(475);
CN_in_sigd(90)	<=	VN_out_sigd(476);
CN_in_sigd(2434)	<=	VN_out_sigd(476);
CN_in_sigd(2698)	<=	VN_out_sigd(476);
CN_in_sigd(4034)	<=	VN_out_sigd(476);
CN_in_sigd(98)	<=	VN_out_sigd(477);
CN_in_sigd(2442)	<=	VN_out_sigd(477);
CN_in_sigd(2706)	<=	VN_out_sigd(477);
CN_in_sigd(4042)	<=	VN_out_sigd(477);
CN_in_sigd(106)	<=	VN_out_sigd(478);
CN_in_sigd(2450)	<=	VN_out_sigd(478);
CN_in_sigd(2714)	<=	VN_out_sigd(478);
CN_in_sigd(4050)	<=	VN_out_sigd(478);
CN_in_sigd(114)	<=	VN_out_sigd(479);
CN_in_sigd(2458)	<=	VN_out_sigd(479);
CN_in_sigd(2722)	<=	VN_out_sigd(479);
CN_in_sigd(4058)	<=	VN_out_sigd(479);
CN_in_sigd(122)	<=	VN_out_sigd(480);
CN_in_sigd(2466)	<=	VN_out_sigd(480);
CN_in_sigd(2730)	<=	VN_out_sigd(480);
CN_in_sigd(4066)	<=	VN_out_sigd(480);
CN_in_sigd(130)	<=	VN_out_sigd(481);
CN_in_sigd(2474)	<=	VN_out_sigd(481);
CN_in_sigd(2738)	<=	VN_out_sigd(481);
CN_in_sigd(4074)	<=	VN_out_sigd(481);
CN_in_sigd(138)	<=	VN_out_sigd(482);
CN_in_sigd(2482)	<=	VN_out_sigd(482);
CN_in_sigd(2746)	<=	VN_out_sigd(482);
CN_in_sigd(4082)	<=	VN_out_sigd(482);
CN_in_sigd(146)	<=	VN_out_sigd(483);
CN_in_sigd(2490)	<=	VN_out_sigd(483);
CN_in_sigd(2754)	<=	VN_out_sigd(483);
CN_in_sigd(4090)	<=	VN_out_sigd(483);
CN_in_sigd(154)	<=	VN_out_sigd(484);
CN_in_sigd(2498)	<=	VN_out_sigd(484);
CN_in_sigd(2762)	<=	VN_out_sigd(484);
CN_in_sigd(4098)	<=	VN_out_sigd(484);
CN_in_sigd(162)	<=	VN_out_sigd(485);
CN_in_sigd(2506)	<=	VN_out_sigd(485);
CN_in_sigd(2770)	<=	VN_out_sigd(485);
CN_in_sigd(4106)	<=	VN_out_sigd(485);
CN_in_sigd(307)	<=	VN_out_sigd(486);
CN_in_sigd(1571)	<=	VN_out_sigd(486);
CN_in_sigd(2875)	<=	VN_out_sigd(486);
CN_in_sigd(4915)	<=	VN_out_sigd(486);
CN_in_sigd(315)	<=	VN_out_sigd(487);
CN_in_sigd(1579)	<=	VN_out_sigd(487);
CN_in_sigd(2883)	<=	VN_out_sigd(487);
CN_in_sigd(4923)	<=	VN_out_sigd(487);
CN_in_sigd(323)	<=	VN_out_sigd(488);
CN_in_sigd(1587)	<=	VN_out_sigd(488);
CN_in_sigd(2891)	<=	VN_out_sigd(488);
CN_in_sigd(4931)	<=	VN_out_sigd(488);
CN_in_sigd(331)	<=	VN_out_sigd(489);
CN_in_sigd(1595)	<=	VN_out_sigd(489);
CN_in_sigd(2899)	<=	VN_out_sigd(489);
CN_in_sigd(4939)	<=	VN_out_sigd(489);
CN_in_sigd(339)	<=	VN_out_sigd(490);
CN_in_sigd(1603)	<=	VN_out_sigd(490);
CN_in_sigd(2907)	<=	VN_out_sigd(490);
CN_in_sigd(4947)	<=	VN_out_sigd(490);
CN_in_sigd(347)	<=	VN_out_sigd(491);
CN_in_sigd(1611)	<=	VN_out_sigd(491);
CN_in_sigd(2915)	<=	VN_out_sigd(491);
CN_in_sigd(4955)	<=	VN_out_sigd(491);
CN_in_sigd(355)	<=	VN_out_sigd(492);
CN_in_sigd(1619)	<=	VN_out_sigd(492);
CN_in_sigd(2923)	<=	VN_out_sigd(492);
CN_in_sigd(4963)	<=	VN_out_sigd(492);
CN_in_sigd(363)	<=	VN_out_sigd(493);
CN_in_sigd(1627)	<=	VN_out_sigd(493);
CN_in_sigd(2931)	<=	VN_out_sigd(493);
CN_in_sigd(4971)	<=	VN_out_sigd(493);
CN_in_sigd(371)	<=	VN_out_sigd(494);
CN_in_sigd(1635)	<=	VN_out_sigd(494);
CN_in_sigd(2939)	<=	VN_out_sigd(494);
CN_in_sigd(4979)	<=	VN_out_sigd(494);
CN_in_sigd(379)	<=	VN_out_sigd(495);
CN_in_sigd(1643)	<=	VN_out_sigd(495);
CN_in_sigd(2947)	<=	VN_out_sigd(495);
CN_in_sigd(4987)	<=	VN_out_sigd(495);
CN_in_sigd(387)	<=	VN_out_sigd(496);
CN_in_sigd(1651)	<=	VN_out_sigd(496);
CN_in_sigd(2955)	<=	VN_out_sigd(496);
CN_in_sigd(4995)	<=	VN_out_sigd(496);
CN_in_sigd(395)	<=	VN_out_sigd(497);
CN_in_sigd(1659)	<=	VN_out_sigd(497);
CN_in_sigd(2963)	<=	VN_out_sigd(497);
CN_in_sigd(5003)	<=	VN_out_sigd(497);
CN_in_sigd(403)	<=	VN_out_sigd(498);
CN_in_sigd(1667)	<=	VN_out_sigd(498);
CN_in_sigd(2971)	<=	VN_out_sigd(498);
CN_in_sigd(5011)	<=	VN_out_sigd(498);
CN_in_sigd(411)	<=	VN_out_sigd(499);
CN_in_sigd(1675)	<=	VN_out_sigd(499);
CN_in_sigd(2979)	<=	VN_out_sigd(499);
CN_in_sigd(5019)	<=	VN_out_sigd(499);
CN_in_sigd(419)	<=	VN_out_sigd(500);
CN_in_sigd(1683)	<=	VN_out_sigd(500);
CN_in_sigd(2987)	<=	VN_out_sigd(500);
CN_in_sigd(5027)	<=	VN_out_sigd(500);
CN_in_sigd(427)	<=	VN_out_sigd(501);
CN_in_sigd(1691)	<=	VN_out_sigd(501);
CN_in_sigd(2995)	<=	VN_out_sigd(501);
CN_in_sigd(5035)	<=	VN_out_sigd(501);
CN_in_sigd(3)	<=	VN_out_sigd(502);
CN_in_sigd(1699)	<=	VN_out_sigd(502);
CN_in_sigd(3003)	<=	VN_out_sigd(502);
CN_in_sigd(5043)	<=	VN_out_sigd(502);
CN_in_sigd(11)	<=	VN_out_sigd(503);
CN_in_sigd(1707)	<=	VN_out_sigd(503);
CN_in_sigd(3011)	<=	VN_out_sigd(503);
CN_in_sigd(5051)	<=	VN_out_sigd(503);
CN_in_sigd(19)	<=	VN_out_sigd(504);
CN_in_sigd(1715)	<=	VN_out_sigd(504);
CN_in_sigd(3019)	<=	VN_out_sigd(504);
CN_in_sigd(5059)	<=	VN_out_sigd(504);
CN_in_sigd(27)	<=	VN_out_sigd(505);
CN_in_sigd(1723)	<=	VN_out_sigd(505);
CN_in_sigd(2595)	<=	VN_out_sigd(505);
CN_in_sigd(5067)	<=	VN_out_sigd(505);
CN_in_sigd(35)	<=	VN_out_sigd(506);
CN_in_sigd(1299)	<=	VN_out_sigd(506);
CN_in_sigd(2603)	<=	VN_out_sigd(506);
CN_in_sigd(5075)	<=	VN_out_sigd(506);
CN_in_sigd(43)	<=	VN_out_sigd(507);
CN_in_sigd(1307)	<=	VN_out_sigd(507);
CN_in_sigd(2611)	<=	VN_out_sigd(507);
CN_in_sigd(5083)	<=	VN_out_sigd(507);
CN_in_sigd(51)	<=	VN_out_sigd(508);
CN_in_sigd(1315)	<=	VN_out_sigd(508);
CN_in_sigd(2619)	<=	VN_out_sigd(508);
CN_in_sigd(5091)	<=	VN_out_sigd(508);
CN_in_sigd(59)	<=	VN_out_sigd(509);
CN_in_sigd(1323)	<=	VN_out_sigd(509);
CN_in_sigd(2627)	<=	VN_out_sigd(509);
CN_in_sigd(5099)	<=	VN_out_sigd(509);
CN_in_sigd(67)	<=	VN_out_sigd(510);
CN_in_sigd(1331)	<=	VN_out_sigd(510);
CN_in_sigd(2635)	<=	VN_out_sigd(510);
CN_in_sigd(5107)	<=	VN_out_sigd(510);
CN_in_sigd(75)	<=	VN_out_sigd(511);
CN_in_sigd(1339)	<=	VN_out_sigd(511);
CN_in_sigd(2643)	<=	VN_out_sigd(511);
CN_in_sigd(5115)	<=	VN_out_sigd(511);
CN_in_sigd(83)	<=	VN_out_sigd(512);
CN_in_sigd(1347)	<=	VN_out_sigd(512);
CN_in_sigd(2651)	<=	VN_out_sigd(512);
CN_in_sigd(5123)	<=	VN_out_sigd(512);
CN_in_sigd(91)	<=	VN_out_sigd(513);
CN_in_sigd(1355)	<=	VN_out_sigd(513);
CN_in_sigd(2659)	<=	VN_out_sigd(513);
CN_in_sigd(5131)	<=	VN_out_sigd(513);
CN_in_sigd(99)	<=	VN_out_sigd(514);
CN_in_sigd(1363)	<=	VN_out_sigd(514);
CN_in_sigd(2667)	<=	VN_out_sigd(514);
CN_in_sigd(5139)	<=	VN_out_sigd(514);
CN_in_sigd(107)	<=	VN_out_sigd(515);
CN_in_sigd(1371)	<=	VN_out_sigd(515);
CN_in_sigd(2675)	<=	VN_out_sigd(515);
CN_in_sigd(5147)	<=	VN_out_sigd(515);
CN_in_sigd(115)	<=	VN_out_sigd(516);
CN_in_sigd(1379)	<=	VN_out_sigd(516);
CN_in_sigd(2683)	<=	VN_out_sigd(516);
CN_in_sigd(5155)	<=	VN_out_sigd(516);
CN_in_sigd(123)	<=	VN_out_sigd(517);
CN_in_sigd(1387)	<=	VN_out_sigd(517);
CN_in_sigd(2691)	<=	VN_out_sigd(517);
CN_in_sigd(5163)	<=	VN_out_sigd(517);
CN_in_sigd(131)	<=	VN_out_sigd(518);
CN_in_sigd(1395)	<=	VN_out_sigd(518);
CN_in_sigd(2699)	<=	VN_out_sigd(518);
CN_in_sigd(5171)	<=	VN_out_sigd(518);
CN_in_sigd(139)	<=	VN_out_sigd(519);
CN_in_sigd(1403)	<=	VN_out_sigd(519);
CN_in_sigd(2707)	<=	VN_out_sigd(519);
CN_in_sigd(5179)	<=	VN_out_sigd(519);
CN_in_sigd(147)	<=	VN_out_sigd(520);
CN_in_sigd(1411)	<=	VN_out_sigd(520);
CN_in_sigd(2715)	<=	VN_out_sigd(520);
CN_in_sigd(4755)	<=	VN_out_sigd(520);
CN_in_sigd(155)	<=	VN_out_sigd(521);
CN_in_sigd(1419)	<=	VN_out_sigd(521);
CN_in_sigd(2723)	<=	VN_out_sigd(521);
CN_in_sigd(4763)	<=	VN_out_sigd(521);
CN_in_sigd(163)	<=	VN_out_sigd(522);
CN_in_sigd(1427)	<=	VN_out_sigd(522);
CN_in_sigd(2731)	<=	VN_out_sigd(522);
CN_in_sigd(4771)	<=	VN_out_sigd(522);
CN_in_sigd(171)	<=	VN_out_sigd(523);
CN_in_sigd(1435)	<=	VN_out_sigd(523);
CN_in_sigd(2739)	<=	VN_out_sigd(523);
CN_in_sigd(4779)	<=	VN_out_sigd(523);
CN_in_sigd(179)	<=	VN_out_sigd(524);
CN_in_sigd(1443)	<=	VN_out_sigd(524);
CN_in_sigd(2747)	<=	VN_out_sigd(524);
CN_in_sigd(4787)	<=	VN_out_sigd(524);
CN_in_sigd(187)	<=	VN_out_sigd(525);
CN_in_sigd(1451)	<=	VN_out_sigd(525);
CN_in_sigd(2755)	<=	VN_out_sigd(525);
CN_in_sigd(4795)	<=	VN_out_sigd(525);
CN_in_sigd(195)	<=	VN_out_sigd(526);
CN_in_sigd(1459)	<=	VN_out_sigd(526);
CN_in_sigd(2763)	<=	VN_out_sigd(526);
CN_in_sigd(4803)	<=	VN_out_sigd(526);
CN_in_sigd(203)	<=	VN_out_sigd(527);
CN_in_sigd(1467)	<=	VN_out_sigd(527);
CN_in_sigd(2771)	<=	VN_out_sigd(527);
CN_in_sigd(4811)	<=	VN_out_sigd(527);
CN_in_sigd(211)	<=	VN_out_sigd(528);
CN_in_sigd(1475)	<=	VN_out_sigd(528);
CN_in_sigd(2779)	<=	VN_out_sigd(528);
CN_in_sigd(4819)	<=	VN_out_sigd(528);
CN_in_sigd(219)	<=	VN_out_sigd(529);
CN_in_sigd(1483)	<=	VN_out_sigd(529);
CN_in_sigd(2787)	<=	VN_out_sigd(529);
CN_in_sigd(4827)	<=	VN_out_sigd(529);
CN_in_sigd(227)	<=	VN_out_sigd(530);
CN_in_sigd(1491)	<=	VN_out_sigd(530);
CN_in_sigd(2795)	<=	VN_out_sigd(530);
CN_in_sigd(4835)	<=	VN_out_sigd(530);
CN_in_sigd(235)	<=	VN_out_sigd(531);
CN_in_sigd(1499)	<=	VN_out_sigd(531);
CN_in_sigd(2803)	<=	VN_out_sigd(531);
CN_in_sigd(4843)	<=	VN_out_sigd(531);
CN_in_sigd(243)	<=	VN_out_sigd(532);
CN_in_sigd(1507)	<=	VN_out_sigd(532);
CN_in_sigd(2811)	<=	VN_out_sigd(532);
CN_in_sigd(4851)	<=	VN_out_sigd(532);
CN_in_sigd(251)	<=	VN_out_sigd(533);
CN_in_sigd(1515)	<=	VN_out_sigd(533);
CN_in_sigd(2819)	<=	VN_out_sigd(533);
CN_in_sigd(4859)	<=	VN_out_sigd(533);
CN_in_sigd(259)	<=	VN_out_sigd(534);
CN_in_sigd(1523)	<=	VN_out_sigd(534);
CN_in_sigd(2827)	<=	VN_out_sigd(534);
CN_in_sigd(4867)	<=	VN_out_sigd(534);
CN_in_sigd(267)	<=	VN_out_sigd(535);
CN_in_sigd(1531)	<=	VN_out_sigd(535);
CN_in_sigd(2835)	<=	VN_out_sigd(535);
CN_in_sigd(4875)	<=	VN_out_sigd(535);
CN_in_sigd(275)	<=	VN_out_sigd(536);
CN_in_sigd(1539)	<=	VN_out_sigd(536);
CN_in_sigd(2843)	<=	VN_out_sigd(536);
CN_in_sigd(4883)	<=	VN_out_sigd(536);
CN_in_sigd(283)	<=	VN_out_sigd(537);
CN_in_sigd(1547)	<=	VN_out_sigd(537);
CN_in_sigd(2851)	<=	VN_out_sigd(537);
CN_in_sigd(4891)	<=	VN_out_sigd(537);
CN_in_sigd(291)	<=	VN_out_sigd(538);
CN_in_sigd(1555)	<=	VN_out_sigd(538);
CN_in_sigd(2859)	<=	VN_out_sigd(538);
CN_in_sigd(4899)	<=	VN_out_sigd(538);
CN_in_sigd(299)	<=	VN_out_sigd(539);
CN_in_sigd(1563)	<=	VN_out_sigd(539);
CN_in_sigd(2867)	<=	VN_out_sigd(539);
CN_in_sigd(4907)	<=	VN_out_sigd(539);
CN_in_sigd(635)	<=	VN_out_sigd(540);
CN_in_sigd(2451)	<=	VN_out_sigd(540);
CN_in_sigd(3419)	<=	VN_out_sigd(540);
CN_in_sigd(4299)	<=	VN_out_sigd(540);
CN_in_sigd(643)	<=	VN_out_sigd(541);
CN_in_sigd(2459)	<=	VN_out_sigd(541);
CN_in_sigd(3427)	<=	VN_out_sigd(541);
CN_in_sigd(4307)	<=	VN_out_sigd(541);
CN_in_sigd(651)	<=	VN_out_sigd(542);
CN_in_sigd(2467)	<=	VN_out_sigd(542);
CN_in_sigd(3435)	<=	VN_out_sigd(542);
CN_in_sigd(4315)	<=	VN_out_sigd(542);
CN_in_sigd(659)	<=	VN_out_sigd(543);
CN_in_sigd(2475)	<=	VN_out_sigd(543);
CN_in_sigd(3443)	<=	VN_out_sigd(543);
CN_in_sigd(3891)	<=	VN_out_sigd(543);
CN_in_sigd(667)	<=	VN_out_sigd(544);
CN_in_sigd(2483)	<=	VN_out_sigd(544);
CN_in_sigd(3451)	<=	VN_out_sigd(544);
CN_in_sigd(3899)	<=	VN_out_sigd(544);
CN_in_sigd(675)	<=	VN_out_sigd(545);
CN_in_sigd(2491)	<=	VN_out_sigd(545);
CN_in_sigd(3027)	<=	VN_out_sigd(545);
CN_in_sigd(3907)	<=	VN_out_sigd(545);
CN_in_sigd(683)	<=	VN_out_sigd(546);
CN_in_sigd(2499)	<=	VN_out_sigd(546);
CN_in_sigd(3035)	<=	VN_out_sigd(546);
CN_in_sigd(3915)	<=	VN_out_sigd(546);
CN_in_sigd(691)	<=	VN_out_sigd(547);
CN_in_sigd(2507)	<=	VN_out_sigd(547);
CN_in_sigd(3043)	<=	VN_out_sigd(547);
CN_in_sigd(3923)	<=	VN_out_sigd(547);
CN_in_sigd(699)	<=	VN_out_sigd(548);
CN_in_sigd(2515)	<=	VN_out_sigd(548);
CN_in_sigd(3051)	<=	VN_out_sigd(548);
CN_in_sigd(3931)	<=	VN_out_sigd(548);
CN_in_sigd(707)	<=	VN_out_sigd(549);
CN_in_sigd(2523)	<=	VN_out_sigd(549);
CN_in_sigd(3059)	<=	VN_out_sigd(549);
CN_in_sigd(3939)	<=	VN_out_sigd(549);
CN_in_sigd(715)	<=	VN_out_sigd(550);
CN_in_sigd(2531)	<=	VN_out_sigd(550);
CN_in_sigd(3067)	<=	VN_out_sigd(550);
CN_in_sigd(3947)	<=	VN_out_sigd(550);
CN_in_sigd(723)	<=	VN_out_sigd(551);
CN_in_sigd(2539)	<=	VN_out_sigd(551);
CN_in_sigd(3075)	<=	VN_out_sigd(551);
CN_in_sigd(3955)	<=	VN_out_sigd(551);
CN_in_sigd(731)	<=	VN_out_sigd(552);
CN_in_sigd(2547)	<=	VN_out_sigd(552);
CN_in_sigd(3083)	<=	VN_out_sigd(552);
CN_in_sigd(3963)	<=	VN_out_sigd(552);
CN_in_sigd(739)	<=	VN_out_sigd(553);
CN_in_sigd(2555)	<=	VN_out_sigd(553);
CN_in_sigd(3091)	<=	VN_out_sigd(553);
CN_in_sigd(3971)	<=	VN_out_sigd(553);
CN_in_sigd(747)	<=	VN_out_sigd(554);
CN_in_sigd(2563)	<=	VN_out_sigd(554);
CN_in_sigd(3099)	<=	VN_out_sigd(554);
CN_in_sigd(3979)	<=	VN_out_sigd(554);
CN_in_sigd(755)	<=	VN_out_sigd(555);
CN_in_sigd(2571)	<=	VN_out_sigd(555);
CN_in_sigd(3107)	<=	VN_out_sigd(555);
CN_in_sigd(3987)	<=	VN_out_sigd(555);
CN_in_sigd(763)	<=	VN_out_sigd(556);
CN_in_sigd(2579)	<=	VN_out_sigd(556);
CN_in_sigd(3115)	<=	VN_out_sigd(556);
CN_in_sigd(3995)	<=	VN_out_sigd(556);
CN_in_sigd(771)	<=	VN_out_sigd(557);
CN_in_sigd(2587)	<=	VN_out_sigd(557);
CN_in_sigd(3123)	<=	VN_out_sigd(557);
CN_in_sigd(4003)	<=	VN_out_sigd(557);
CN_in_sigd(779)	<=	VN_out_sigd(558);
CN_in_sigd(2163)	<=	VN_out_sigd(558);
CN_in_sigd(3131)	<=	VN_out_sigd(558);
CN_in_sigd(4011)	<=	VN_out_sigd(558);
CN_in_sigd(787)	<=	VN_out_sigd(559);
CN_in_sigd(2171)	<=	VN_out_sigd(559);
CN_in_sigd(3139)	<=	VN_out_sigd(559);
CN_in_sigd(4019)	<=	VN_out_sigd(559);
CN_in_sigd(795)	<=	VN_out_sigd(560);
CN_in_sigd(2179)	<=	VN_out_sigd(560);
CN_in_sigd(3147)	<=	VN_out_sigd(560);
CN_in_sigd(4027)	<=	VN_out_sigd(560);
CN_in_sigd(803)	<=	VN_out_sigd(561);
CN_in_sigd(2187)	<=	VN_out_sigd(561);
CN_in_sigd(3155)	<=	VN_out_sigd(561);
CN_in_sigd(4035)	<=	VN_out_sigd(561);
CN_in_sigd(811)	<=	VN_out_sigd(562);
CN_in_sigd(2195)	<=	VN_out_sigd(562);
CN_in_sigd(3163)	<=	VN_out_sigd(562);
CN_in_sigd(4043)	<=	VN_out_sigd(562);
CN_in_sigd(819)	<=	VN_out_sigd(563);
CN_in_sigd(2203)	<=	VN_out_sigd(563);
CN_in_sigd(3171)	<=	VN_out_sigd(563);
CN_in_sigd(4051)	<=	VN_out_sigd(563);
CN_in_sigd(827)	<=	VN_out_sigd(564);
CN_in_sigd(2211)	<=	VN_out_sigd(564);
CN_in_sigd(3179)	<=	VN_out_sigd(564);
CN_in_sigd(4059)	<=	VN_out_sigd(564);
CN_in_sigd(835)	<=	VN_out_sigd(565);
CN_in_sigd(2219)	<=	VN_out_sigd(565);
CN_in_sigd(3187)	<=	VN_out_sigd(565);
CN_in_sigd(4067)	<=	VN_out_sigd(565);
CN_in_sigd(843)	<=	VN_out_sigd(566);
CN_in_sigd(2227)	<=	VN_out_sigd(566);
CN_in_sigd(3195)	<=	VN_out_sigd(566);
CN_in_sigd(4075)	<=	VN_out_sigd(566);
CN_in_sigd(851)	<=	VN_out_sigd(567);
CN_in_sigd(2235)	<=	VN_out_sigd(567);
CN_in_sigd(3203)	<=	VN_out_sigd(567);
CN_in_sigd(4083)	<=	VN_out_sigd(567);
CN_in_sigd(859)	<=	VN_out_sigd(568);
CN_in_sigd(2243)	<=	VN_out_sigd(568);
CN_in_sigd(3211)	<=	VN_out_sigd(568);
CN_in_sigd(4091)	<=	VN_out_sigd(568);
CN_in_sigd(435)	<=	VN_out_sigd(569);
CN_in_sigd(2251)	<=	VN_out_sigd(569);
CN_in_sigd(3219)	<=	VN_out_sigd(569);
CN_in_sigd(4099)	<=	VN_out_sigd(569);
CN_in_sigd(443)	<=	VN_out_sigd(570);
CN_in_sigd(2259)	<=	VN_out_sigd(570);
CN_in_sigd(3227)	<=	VN_out_sigd(570);
CN_in_sigd(4107)	<=	VN_out_sigd(570);
CN_in_sigd(451)	<=	VN_out_sigd(571);
CN_in_sigd(2267)	<=	VN_out_sigd(571);
CN_in_sigd(3235)	<=	VN_out_sigd(571);
CN_in_sigd(4115)	<=	VN_out_sigd(571);
CN_in_sigd(459)	<=	VN_out_sigd(572);
CN_in_sigd(2275)	<=	VN_out_sigd(572);
CN_in_sigd(3243)	<=	VN_out_sigd(572);
CN_in_sigd(4123)	<=	VN_out_sigd(572);
CN_in_sigd(467)	<=	VN_out_sigd(573);
CN_in_sigd(2283)	<=	VN_out_sigd(573);
CN_in_sigd(3251)	<=	VN_out_sigd(573);
CN_in_sigd(4131)	<=	VN_out_sigd(573);
CN_in_sigd(475)	<=	VN_out_sigd(574);
CN_in_sigd(2291)	<=	VN_out_sigd(574);
CN_in_sigd(3259)	<=	VN_out_sigd(574);
CN_in_sigd(4139)	<=	VN_out_sigd(574);
CN_in_sigd(483)	<=	VN_out_sigd(575);
CN_in_sigd(2299)	<=	VN_out_sigd(575);
CN_in_sigd(3267)	<=	VN_out_sigd(575);
CN_in_sigd(4147)	<=	VN_out_sigd(575);
CN_in_sigd(491)	<=	VN_out_sigd(576);
CN_in_sigd(2307)	<=	VN_out_sigd(576);
CN_in_sigd(3275)	<=	VN_out_sigd(576);
CN_in_sigd(4155)	<=	VN_out_sigd(576);
CN_in_sigd(499)	<=	VN_out_sigd(577);
CN_in_sigd(2315)	<=	VN_out_sigd(577);
CN_in_sigd(3283)	<=	VN_out_sigd(577);
CN_in_sigd(4163)	<=	VN_out_sigd(577);
CN_in_sigd(507)	<=	VN_out_sigd(578);
CN_in_sigd(2323)	<=	VN_out_sigd(578);
CN_in_sigd(3291)	<=	VN_out_sigd(578);
CN_in_sigd(4171)	<=	VN_out_sigd(578);
CN_in_sigd(515)	<=	VN_out_sigd(579);
CN_in_sigd(2331)	<=	VN_out_sigd(579);
CN_in_sigd(3299)	<=	VN_out_sigd(579);
CN_in_sigd(4179)	<=	VN_out_sigd(579);
CN_in_sigd(523)	<=	VN_out_sigd(580);
CN_in_sigd(2339)	<=	VN_out_sigd(580);
CN_in_sigd(3307)	<=	VN_out_sigd(580);
CN_in_sigd(4187)	<=	VN_out_sigd(580);
CN_in_sigd(531)	<=	VN_out_sigd(581);
CN_in_sigd(2347)	<=	VN_out_sigd(581);
CN_in_sigd(3315)	<=	VN_out_sigd(581);
CN_in_sigd(4195)	<=	VN_out_sigd(581);
CN_in_sigd(539)	<=	VN_out_sigd(582);
CN_in_sigd(2355)	<=	VN_out_sigd(582);
CN_in_sigd(3323)	<=	VN_out_sigd(582);
CN_in_sigd(4203)	<=	VN_out_sigd(582);
CN_in_sigd(547)	<=	VN_out_sigd(583);
CN_in_sigd(2363)	<=	VN_out_sigd(583);
CN_in_sigd(3331)	<=	VN_out_sigd(583);
CN_in_sigd(4211)	<=	VN_out_sigd(583);
CN_in_sigd(555)	<=	VN_out_sigd(584);
CN_in_sigd(2371)	<=	VN_out_sigd(584);
CN_in_sigd(3339)	<=	VN_out_sigd(584);
CN_in_sigd(4219)	<=	VN_out_sigd(584);
CN_in_sigd(563)	<=	VN_out_sigd(585);
CN_in_sigd(2379)	<=	VN_out_sigd(585);
CN_in_sigd(3347)	<=	VN_out_sigd(585);
CN_in_sigd(4227)	<=	VN_out_sigd(585);
CN_in_sigd(571)	<=	VN_out_sigd(586);
CN_in_sigd(2387)	<=	VN_out_sigd(586);
CN_in_sigd(3355)	<=	VN_out_sigd(586);
CN_in_sigd(4235)	<=	VN_out_sigd(586);
CN_in_sigd(579)	<=	VN_out_sigd(587);
CN_in_sigd(2395)	<=	VN_out_sigd(587);
CN_in_sigd(3363)	<=	VN_out_sigd(587);
CN_in_sigd(4243)	<=	VN_out_sigd(587);
CN_in_sigd(587)	<=	VN_out_sigd(588);
CN_in_sigd(2403)	<=	VN_out_sigd(588);
CN_in_sigd(3371)	<=	VN_out_sigd(588);
CN_in_sigd(4251)	<=	VN_out_sigd(588);
CN_in_sigd(595)	<=	VN_out_sigd(589);
CN_in_sigd(2411)	<=	VN_out_sigd(589);
CN_in_sigd(3379)	<=	VN_out_sigd(589);
CN_in_sigd(4259)	<=	VN_out_sigd(589);
CN_in_sigd(603)	<=	VN_out_sigd(590);
CN_in_sigd(2419)	<=	VN_out_sigd(590);
CN_in_sigd(3387)	<=	VN_out_sigd(590);
CN_in_sigd(4267)	<=	VN_out_sigd(590);
CN_in_sigd(611)	<=	VN_out_sigd(591);
CN_in_sigd(2427)	<=	VN_out_sigd(591);
CN_in_sigd(3395)	<=	VN_out_sigd(591);
CN_in_sigd(4275)	<=	VN_out_sigd(591);
CN_in_sigd(619)	<=	VN_out_sigd(592);
CN_in_sigd(2435)	<=	VN_out_sigd(592);
CN_in_sigd(3403)	<=	VN_out_sigd(592);
CN_in_sigd(4283)	<=	VN_out_sigd(592);
CN_in_sigd(627)	<=	VN_out_sigd(593);
CN_in_sigd(2443)	<=	VN_out_sigd(593);
CN_in_sigd(3411)	<=	VN_out_sigd(593);
CN_in_sigd(4291)	<=	VN_out_sigd(593);
CN_in_sigd(1283)	<=	VN_out_sigd(594);
CN_in_sigd(1811)	<=	VN_out_sigd(594);
CN_in_sigd(3883)	<=	VN_out_sigd(594);
CN_in_sigd(4651)	<=	VN_out_sigd(594);
CN_in_sigd(1291)	<=	VN_out_sigd(595);
CN_in_sigd(1819)	<=	VN_out_sigd(595);
CN_in_sigd(3459)	<=	VN_out_sigd(595);
CN_in_sigd(4659)	<=	VN_out_sigd(595);
CN_in_sigd(867)	<=	VN_out_sigd(596);
CN_in_sigd(1827)	<=	VN_out_sigd(596);
CN_in_sigd(3467)	<=	VN_out_sigd(596);
CN_in_sigd(4667)	<=	VN_out_sigd(596);
CN_in_sigd(875)	<=	VN_out_sigd(597);
CN_in_sigd(1835)	<=	VN_out_sigd(597);
CN_in_sigd(3475)	<=	VN_out_sigd(597);
CN_in_sigd(4675)	<=	VN_out_sigd(597);
CN_in_sigd(883)	<=	VN_out_sigd(598);
CN_in_sigd(1843)	<=	VN_out_sigd(598);
CN_in_sigd(3483)	<=	VN_out_sigd(598);
CN_in_sigd(4683)	<=	VN_out_sigd(598);
CN_in_sigd(891)	<=	VN_out_sigd(599);
CN_in_sigd(1851)	<=	VN_out_sigd(599);
CN_in_sigd(3491)	<=	VN_out_sigd(599);
CN_in_sigd(4691)	<=	VN_out_sigd(599);
CN_in_sigd(899)	<=	VN_out_sigd(600);
CN_in_sigd(1859)	<=	VN_out_sigd(600);
CN_in_sigd(3499)	<=	VN_out_sigd(600);
CN_in_sigd(4699)	<=	VN_out_sigd(600);
CN_in_sigd(907)	<=	VN_out_sigd(601);
CN_in_sigd(1867)	<=	VN_out_sigd(601);
CN_in_sigd(3507)	<=	VN_out_sigd(601);
CN_in_sigd(4707)	<=	VN_out_sigd(601);
CN_in_sigd(915)	<=	VN_out_sigd(602);
CN_in_sigd(1875)	<=	VN_out_sigd(602);
CN_in_sigd(3515)	<=	VN_out_sigd(602);
CN_in_sigd(4715)	<=	VN_out_sigd(602);
CN_in_sigd(923)	<=	VN_out_sigd(603);
CN_in_sigd(1883)	<=	VN_out_sigd(603);
CN_in_sigd(3523)	<=	VN_out_sigd(603);
CN_in_sigd(4723)	<=	VN_out_sigd(603);
CN_in_sigd(931)	<=	VN_out_sigd(604);
CN_in_sigd(1891)	<=	VN_out_sigd(604);
CN_in_sigd(3531)	<=	VN_out_sigd(604);
CN_in_sigd(4731)	<=	VN_out_sigd(604);
CN_in_sigd(939)	<=	VN_out_sigd(605);
CN_in_sigd(1899)	<=	VN_out_sigd(605);
CN_in_sigd(3539)	<=	VN_out_sigd(605);
CN_in_sigd(4739)	<=	VN_out_sigd(605);
CN_in_sigd(947)	<=	VN_out_sigd(606);
CN_in_sigd(1907)	<=	VN_out_sigd(606);
CN_in_sigd(3547)	<=	VN_out_sigd(606);
CN_in_sigd(4747)	<=	VN_out_sigd(606);
CN_in_sigd(955)	<=	VN_out_sigd(607);
CN_in_sigd(1915)	<=	VN_out_sigd(607);
CN_in_sigd(3555)	<=	VN_out_sigd(607);
CN_in_sigd(4323)	<=	VN_out_sigd(607);
CN_in_sigd(963)	<=	VN_out_sigd(608);
CN_in_sigd(1923)	<=	VN_out_sigd(608);
CN_in_sigd(3563)	<=	VN_out_sigd(608);
CN_in_sigd(4331)	<=	VN_out_sigd(608);
CN_in_sigd(971)	<=	VN_out_sigd(609);
CN_in_sigd(1931)	<=	VN_out_sigd(609);
CN_in_sigd(3571)	<=	VN_out_sigd(609);
CN_in_sigd(4339)	<=	VN_out_sigd(609);
CN_in_sigd(979)	<=	VN_out_sigd(610);
CN_in_sigd(1939)	<=	VN_out_sigd(610);
CN_in_sigd(3579)	<=	VN_out_sigd(610);
CN_in_sigd(4347)	<=	VN_out_sigd(610);
CN_in_sigd(987)	<=	VN_out_sigd(611);
CN_in_sigd(1947)	<=	VN_out_sigd(611);
CN_in_sigd(3587)	<=	VN_out_sigd(611);
CN_in_sigd(4355)	<=	VN_out_sigd(611);
CN_in_sigd(995)	<=	VN_out_sigd(612);
CN_in_sigd(1955)	<=	VN_out_sigd(612);
CN_in_sigd(3595)	<=	VN_out_sigd(612);
CN_in_sigd(4363)	<=	VN_out_sigd(612);
CN_in_sigd(1003)	<=	VN_out_sigd(613);
CN_in_sigd(1963)	<=	VN_out_sigd(613);
CN_in_sigd(3603)	<=	VN_out_sigd(613);
CN_in_sigd(4371)	<=	VN_out_sigd(613);
CN_in_sigd(1011)	<=	VN_out_sigd(614);
CN_in_sigd(1971)	<=	VN_out_sigd(614);
CN_in_sigd(3611)	<=	VN_out_sigd(614);
CN_in_sigd(4379)	<=	VN_out_sigd(614);
CN_in_sigd(1019)	<=	VN_out_sigd(615);
CN_in_sigd(1979)	<=	VN_out_sigd(615);
CN_in_sigd(3619)	<=	VN_out_sigd(615);
CN_in_sigd(4387)	<=	VN_out_sigd(615);
CN_in_sigd(1027)	<=	VN_out_sigd(616);
CN_in_sigd(1987)	<=	VN_out_sigd(616);
CN_in_sigd(3627)	<=	VN_out_sigd(616);
CN_in_sigd(4395)	<=	VN_out_sigd(616);
CN_in_sigd(1035)	<=	VN_out_sigd(617);
CN_in_sigd(1995)	<=	VN_out_sigd(617);
CN_in_sigd(3635)	<=	VN_out_sigd(617);
CN_in_sigd(4403)	<=	VN_out_sigd(617);
CN_in_sigd(1043)	<=	VN_out_sigd(618);
CN_in_sigd(2003)	<=	VN_out_sigd(618);
CN_in_sigd(3643)	<=	VN_out_sigd(618);
CN_in_sigd(4411)	<=	VN_out_sigd(618);
CN_in_sigd(1051)	<=	VN_out_sigd(619);
CN_in_sigd(2011)	<=	VN_out_sigd(619);
CN_in_sigd(3651)	<=	VN_out_sigd(619);
CN_in_sigd(4419)	<=	VN_out_sigd(619);
CN_in_sigd(1059)	<=	VN_out_sigd(620);
CN_in_sigd(2019)	<=	VN_out_sigd(620);
CN_in_sigd(3659)	<=	VN_out_sigd(620);
CN_in_sigd(4427)	<=	VN_out_sigd(620);
CN_in_sigd(1067)	<=	VN_out_sigd(621);
CN_in_sigd(2027)	<=	VN_out_sigd(621);
CN_in_sigd(3667)	<=	VN_out_sigd(621);
CN_in_sigd(4435)	<=	VN_out_sigd(621);
CN_in_sigd(1075)	<=	VN_out_sigd(622);
CN_in_sigd(2035)	<=	VN_out_sigd(622);
CN_in_sigd(3675)	<=	VN_out_sigd(622);
CN_in_sigd(4443)	<=	VN_out_sigd(622);
CN_in_sigd(1083)	<=	VN_out_sigd(623);
CN_in_sigd(2043)	<=	VN_out_sigd(623);
CN_in_sigd(3683)	<=	VN_out_sigd(623);
CN_in_sigd(4451)	<=	VN_out_sigd(623);
CN_in_sigd(1091)	<=	VN_out_sigd(624);
CN_in_sigd(2051)	<=	VN_out_sigd(624);
CN_in_sigd(3691)	<=	VN_out_sigd(624);
CN_in_sigd(4459)	<=	VN_out_sigd(624);
CN_in_sigd(1099)	<=	VN_out_sigd(625);
CN_in_sigd(2059)	<=	VN_out_sigd(625);
CN_in_sigd(3699)	<=	VN_out_sigd(625);
CN_in_sigd(4467)	<=	VN_out_sigd(625);
CN_in_sigd(1107)	<=	VN_out_sigd(626);
CN_in_sigd(2067)	<=	VN_out_sigd(626);
CN_in_sigd(3707)	<=	VN_out_sigd(626);
CN_in_sigd(4475)	<=	VN_out_sigd(626);
CN_in_sigd(1115)	<=	VN_out_sigd(627);
CN_in_sigd(2075)	<=	VN_out_sigd(627);
CN_in_sigd(3715)	<=	VN_out_sigd(627);
CN_in_sigd(4483)	<=	VN_out_sigd(627);
CN_in_sigd(1123)	<=	VN_out_sigd(628);
CN_in_sigd(2083)	<=	VN_out_sigd(628);
CN_in_sigd(3723)	<=	VN_out_sigd(628);
CN_in_sigd(4491)	<=	VN_out_sigd(628);
CN_in_sigd(1131)	<=	VN_out_sigd(629);
CN_in_sigd(2091)	<=	VN_out_sigd(629);
CN_in_sigd(3731)	<=	VN_out_sigd(629);
CN_in_sigd(4499)	<=	VN_out_sigd(629);
CN_in_sigd(1139)	<=	VN_out_sigd(630);
CN_in_sigd(2099)	<=	VN_out_sigd(630);
CN_in_sigd(3739)	<=	VN_out_sigd(630);
CN_in_sigd(4507)	<=	VN_out_sigd(630);
CN_in_sigd(1147)	<=	VN_out_sigd(631);
CN_in_sigd(2107)	<=	VN_out_sigd(631);
CN_in_sigd(3747)	<=	VN_out_sigd(631);
CN_in_sigd(4515)	<=	VN_out_sigd(631);
CN_in_sigd(1155)	<=	VN_out_sigd(632);
CN_in_sigd(2115)	<=	VN_out_sigd(632);
CN_in_sigd(3755)	<=	VN_out_sigd(632);
CN_in_sigd(4523)	<=	VN_out_sigd(632);
CN_in_sigd(1163)	<=	VN_out_sigd(633);
CN_in_sigd(2123)	<=	VN_out_sigd(633);
CN_in_sigd(3763)	<=	VN_out_sigd(633);
CN_in_sigd(4531)	<=	VN_out_sigd(633);
CN_in_sigd(1171)	<=	VN_out_sigd(634);
CN_in_sigd(2131)	<=	VN_out_sigd(634);
CN_in_sigd(3771)	<=	VN_out_sigd(634);
CN_in_sigd(4539)	<=	VN_out_sigd(634);
CN_in_sigd(1179)	<=	VN_out_sigd(635);
CN_in_sigd(2139)	<=	VN_out_sigd(635);
CN_in_sigd(3779)	<=	VN_out_sigd(635);
CN_in_sigd(4547)	<=	VN_out_sigd(635);
CN_in_sigd(1187)	<=	VN_out_sigd(636);
CN_in_sigd(2147)	<=	VN_out_sigd(636);
CN_in_sigd(3787)	<=	VN_out_sigd(636);
CN_in_sigd(4555)	<=	VN_out_sigd(636);
CN_in_sigd(1195)	<=	VN_out_sigd(637);
CN_in_sigd(2155)	<=	VN_out_sigd(637);
CN_in_sigd(3795)	<=	VN_out_sigd(637);
CN_in_sigd(4563)	<=	VN_out_sigd(637);
CN_in_sigd(1203)	<=	VN_out_sigd(638);
CN_in_sigd(1731)	<=	VN_out_sigd(638);
CN_in_sigd(3803)	<=	VN_out_sigd(638);
CN_in_sigd(4571)	<=	VN_out_sigd(638);
CN_in_sigd(1211)	<=	VN_out_sigd(639);
CN_in_sigd(1739)	<=	VN_out_sigd(639);
CN_in_sigd(3811)	<=	VN_out_sigd(639);
CN_in_sigd(4579)	<=	VN_out_sigd(639);
CN_in_sigd(1219)	<=	VN_out_sigd(640);
CN_in_sigd(1747)	<=	VN_out_sigd(640);
CN_in_sigd(3819)	<=	VN_out_sigd(640);
CN_in_sigd(4587)	<=	VN_out_sigd(640);
CN_in_sigd(1227)	<=	VN_out_sigd(641);
CN_in_sigd(1755)	<=	VN_out_sigd(641);
CN_in_sigd(3827)	<=	VN_out_sigd(641);
CN_in_sigd(4595)	<=	VN_out_sigd(641);
CN_in_sigd(1235)	<=	VN_out_sigd(642);
CN_in_sigd(1763)	<=	VN_out_sigd(642);
CN_in_sigd(3835)	<=	VN_out_sigd(642);
CN_in_sigd(4603)	<=	VN_out_sigd(642);
CN_in_sigd(1243)	<=	VN_out_sigd(643);
CN_in_sigd(1771)	<=	VN_out_sigd(643);
CN_in_sigd(3843)	<=	VN_out_sigd(643);
CN_in_sigd(4611)	<=	VN_out_sigd(643);
CN_in_sigd(1251)	<=	VN_out_sigd(644);
CN_in_sigd(1779)	<=	VN_out_sigd(644);
CN_in_sigd(3851)	<=	VN_out_sigd(644);
CN_in_sigd(4619)	<=	VN_out_sigd(644);
CN_in_sigd(1259)	<=	VN_out_sigd(645);
CN_in_sigd(1787)	<=	VN_out_sigd(645);
CN_in_sigd(3859)	<=	VN_out_sigd(645);
CN_in_sigd(4627)	<=	VN_out_sigd(645);
CN_in_sigd(1267)	<=	VN_out_sigd(646);
CN_in_sigd(1795)	<=	VN_out_sigd(646);
CN_in_sigd(3867)	<=	VN_out_sigd(646);
CN_in_sigd(4635)	<=	VN_out_sigd(646);
CN_in_sigd(1275)	<=	VN_out_sigd(647);
CN_in_sigd(1803)	<=	VN_out_sigd(647);
CN_in_sigd(3875)	<=	VN_out_sigd(647);
CN_in_sigd(4643)	<=	VN_out_sigd(647);
CN_in_sigd(900)	<=	VN_out_sigd(648);
CN_in_sigd(2580)	<=	VN_out_sigd(648);
CN_in_sigd(3004)	<=	VN_out_sigd(648);
CN_in_sigd(4420)	<=	VN_out_sigd(648);
CN_in_sigd(908)	<=	VN_out_sigd(649);
CN_in_sigd(2588)	<=	VN_out_sigd(649);
CN_in_sigd(3012)	<=	VN_out_sigd(649);
CN_in_sigd(4428)	<=	VN_out_sigd(649);
CN_in_sigd(916)	<=	VN_out_sigd(650);
CN_in_sigd(2164)	<=	VN_out_sigd(650);
CN_in_sigd(3020)	<=	VN_out_sigd(650);
CN_in_sigd(4436)	<=	VN_out_sigd(650);
CN_in_sigd(924)	<=	VN_out_sigd(651);
CN_in_sigd(2172)	<=	VN_out_sigd(651);
CN_in_sigd(2596)	<=	VN_out_sigd(651);
CN_in_sigd(4444)	<=	VN_out_sigd(651);
CN_in_sigd(932)	<=	VN_out_sigd(652);
CN_in_sigd(2180)	<=	VN_out_sigd(652);
CN_in_sigd(2604)	<=	VN_out_sigd(652);
CN_in_sigd(4452)	<=	VN_out_sigd(652);
CN_in_sigd(940)	<=	VN_out_sigd(653);
CN_in_sigd(2188)	<=	VN_out_sigd(653);
CN_in_sigd(2612)	<=	VN_out_sigd(653);
CN_in_sigd(4460)	<=	VN_out_sigd(653);
CN_in_sigd(948)	<=	VN_out_sigd(654);
CN_in_sigd(2196)	<=	VN_out_sigd(654);
CN_in_sigd(2620)	<=	VN_out_sigd(654);
CN_in_sigd(4468)	<=	VN_out_sigd(654);
CN_in_sigd(956)	<=	VN_out_sigd(655);
CN_in_sigd(2204)	<=	VN_out_sigd(655);
CN_in_sigd(2628)	<=	VN_out_sigd(655);
CN_in_sigd(4476)	<=	VN_out_sigd(655);
CN_in_sigd(964)	<=	VN_out_sigd(656);
CN_in_sigd(2212)	<=	VN_out_sigd(656);
CN_in_sigd(2636)	<=	VN_out_sigd(656);
CN_in_sigd(4484)	<=	VN_out_sigd(656);
CN_in_sigd(972)	<=	VN_out_sigd(657);
CN_in_sigd(2220)	<=	VN_out_sigd(657);
CN_in_sigd(2644)	<=	VN_out_sigd(657);
CN_in_sigd(4492)	<=	VN_out_sigd(657);
CN_in_sigd(980)	<=	VN_out_sigd(658);
CN_in_sigd(2228)	<=	VN_out_sigd(658);
CN_in_sigd(2652)	<=	VN_out_sigd(658);
CN_in_sigd(4500)	<=	VN_out_sigd(658);
CN_in_sigd(988)	<=	VN_out_sigd(659);
CN_in_sigd(2236)	<=	VN_out_sigd(659);
CN_in_sigd(2660)	<=	VN_out_sigd(659);
CN_in_sigd(4508)	<=	VN_out_sigd(659);
CN_in_sigd(996)	<=	VN_out_sigd(660);
CN_in_sigd(2244)	<=	VN_out_sigd(660);
CN_in_sigd(2668)	<=	VN_out_sigd(660);
CN_in_sigd(4516)	<=	VN_out_sigd(660);
CN_in_sigd(1004)	<=	VN_out_sigd(661);
CN_in_sigd(2252)	<=	VN_out_sigd(661);
CN_in_sigd(2676)	<=	VN_out_sigd(661);
CN_in_sigd(4524)	<=	VN_out_sigd(661);
CN_in_sigd(1012)	<=	VN_out_sigd(662);
CN_in_sigd(2260)	<=	VN_out_sigd(662);
CN_in_sigd(2684)	<=	VN_out_sigd(662);
CN_in_sigd(4532)	<=	VN_out_sigd(662);
CN_in_sigd(1020)	<=	VN_out_sigd(663);
CN_in_sigd(2268)	<=	VN_out_sigd(663);
CN_in_sigd(2692)	<=	VN_out_sigd(663);
CN_in_sigd(4540)	<=	VN_out_sigd(663);
CN_in_sigd(1028)	<=	VN_out_sigd(664);
CN_in_sigd(2276)	<=	VN_out_sigd(664);
CN_in_sigd(2700)	<=	VN_out_sigd(664);
CN_in_sigd(4548)	<=	VN_out_sigd(664);
CN_in_sigd(1036)	<=	VN_out_sigd(665);
CN_in_sigd(2284)	<=	VN_out_sigd(665);
CN_in_sigd(2708)	<=	VN_out_sigd(665);
CN_in_sigd(4556)	<=	VN_out_sigd(665);
CN_in_sigd(1044)	<=	VN_out_sigd(666);
CN_in_sigd(2292)	<=	VN_out_sigd(666);
CN_in_sigd(2716)	<=	VN_out_sigd(666);
CN_in_sigd(4564)	<=	VN_out_sigd(666);
CN_in_sigd(1052)	<=	VN_out_sigd(667);
CN_in_sigd(2300)	<=	VN_out_sigd(667);
CN_in_sigd(2724)	<=	VN_out_sigd(667);
CN_in_sigd(4572)	<=	VN_out_sigd(667);
CN_in_sigd(1060)	<=	VN_out_sigd(668);
CN_in_sigd(2308)	<=	VN_out_sigd(668);
CN_in_sigd(2732)	<=	VN_out_sigd(668);
CN_in_sigd(4580)	<=	VN_out_sigd(668);
CN_in_sigd(1068)	<=	VN_out_sigd(669);
CN_in_sigd(2316)	<=	VN_out_sigd(669);
CN_in_sigd(2740)	<=	VN_out_sigd(669);
CN_in_sigd(4588)	<=	VN_out_sigd(669);
CN_in_sigd(1076)	<=	VN_out_sigd(670);
CN_in_sigd(2324)	<=	VN_out_sigd(670);
CN_in_sigd(2748)	<=	VN_out_sigd(670);
CN_in_sigd(4596)	<=	VN_out_sigd(670);
CN_in_sigd(1084)	<=	VN_out_sigd(671);
CN_in_sigd(2332)	<=	VN_out_sigd(671);
CN_in_sigd(2756)	<=	VN_out_sigd(671);
CN_in_sigd(4604)	<=	VN_out_sigd(671);
CN_in_sigd(1092)	<=	VN_out_sigd(672);
CN_in_sigd(2340)	<=	VN_out_sigd(672);
CN_in_sigd(2764)	<=	VN_out_sigd(672);
CN_in_sigd(4612)	<=	VN_out_sigd(672);
CN_in_sigd(1100)	<=	VN_out_sigd(673);
CN_in_sigd(2348)	<=	VN_out_sigd(673);
CN_in_sigd(2772)	<=	VN_out_sigd(673);
CN_in_sigd(4620)	<=	VN_out_sigd(673);
CN_in_sigd(1108)	<=	VN_out_sigd(674);
CN_in_sigd(2356)	<=	VN_out_sigd(674);
CN_in_sigd(2780)	<=	VN_out_sigd(674);
CN_in_sigd(4628)	<=	VN_out_sigd(674);
CN_in_sigd(1116)	<=	VN_out_sigd(675);
CN_in_sigd(2364)	<=	VN_out_sigd(675);
CN_in_sigd(2788)	<=	VN_out_sigd(675);
CN_in_sigd(4636)	<=	VN_out_sigd(675);
CN_in_sigd(1124)	<=	VN_out_sigd(676);
CN_in_sigd(2372)	<=	VN_out_sigd(676);
CN_in_sigd(2796)	<=	VN_out_sigd(676);
CN_in_sigd(4644)	<=	VN_out_sigd(676);
CN_in_sigd(1132)	<=	VN_out_sigd(677);
CN_in_sigd(2380)	<=	VN_out_sigd(677);
CN_in_sigd(2804)	<=	VN_out_sigd(677);
CN_in_sigd(4652)	<=	VN_out_sigd(677);
CN_in_sigd(1140)	<=	VN_out_sigd(678);
CN_in_sigd(2388)	<=	VN_out_sigd(678);
CN_in_sigd(2812)	<=	VN_out_sigd(678);
CN_in_sigd(4660)	<=	VN_out_sigd(678);
CN_in_sigd(1148)	<=	VN_out_sigd(679);
CN_in_sigd(2396)	<=	VN_out_sigd(679);
CN_in_sigd(2820)	<=	VN_out_sigd(679);
CN_in_sigd(4668)	<=	VN_out_sigd(679);
CN_in_sigd(1156)	<=	VN_out_sigd(680);
CN_in_sigd(2404)	<=	VN_out_sigd(680);
CN_in_sigd(2828)	<=	VN_out_sigd(680);
CN_in_sigd(4676)	<=	VN_out_sigd(680);
CN_in_sigd(1164)	<=	VN_out_sigd(681);
CN_in_sigd(2412)	<=	VN_out_sigd(681);
CN_in_sigd(2836)	<=	VN_out_sigd(681);
CN_in_sigd(4684)	<=	VN_out_sigd(681);
CN_in_sigd(1172)	<=	VN_out_sigd(682);
CN_in_sigd(2420)	<=	VN_out_sigd(682);
CN_in_sigd(2844)	<=	VN_out_sigd(682);
CN_in_sigd(4692)	<=	VN_out_sigd(682);
CN_in_sigd(1180)	<=	VN_out_sigd(683);
CN_in_sigd(2428)	<=	VN_out_sigd(683);
CN_in_sigd(2852)	<=	VN_out_sigd(683);
CN_in_sigd(4700)	<=	VN_out_sigd(683);
CN_in_sigd(1188)	<=	VN_out_sigd(684);
CN_in_sigd(2436)	<=	VN_out_sigd(684);
CN_in_sigd(2860)	<=	VN_out_sigd(684);
CN_in_sigd(4708)	<=	VN_out_sigd(684);
CN_in_sigd(1196)	<=	VN_out_sigd(685);
CN_in_sigd(2444)	<=	VN_out_sigd(685);
CN_in_sigd(2868)	<=	VN_out_sigd(685);
CN_in_sigd(4716)	<=	VN_out_sigd(685);
CN_in_sigd(1204)	<=	VN_out_sigd(686);
CN_in_sigd(2452)	<=	VN_out_sigd(686);
CN_in_sigd(2876)	<=	VN_out_sigd(686);
CN_in_sigd(4724)	<=	VN_out_sigd(686);
CN_in_sigd(1212)	<=	VN_out_sigd(687);
CN_in_sigd(2460)	<=	VN_out_sigd(687);
CN_in_sigd(2884)	<=	VN_out_sigd(687);
CN_in_sigd(4732)	<=	VN_out_sigd(687);
CN_in_sigd(1220)	<=	VN_out_sigd(688);
CN_in_sigd(2468)	<=	VN_out_sigd(688);
CN_in_sigd(2892)	<=	VN_out_sigd(688);
CN_in_sigd(4740)	<=	VN_out_sigd(688);
CN_in_sigd(1228)	<=	VN_out_sigd(689);
CN_in_sigd(2476)	<=	VN_out_sigd(689);
CN_in_sigd(2900)	<=	VN_out_sigd(689);
CN_in_sigd(4748)	<=	VN_out_sigd(689);
CN_in_sigd(1236)	<=	VN_out_sigd(690);
CN_in_sigd(2484)	<=	VN_out_sigd(690);
CN_in_sigd(2908)	<=	VN_out_sigd(690);
CN_in_sigd(4324)	<=	VN_out_sigd(690);
CN_in_sigd(1244)	<=	VN_out_sigd(691);
CN_in_sigd(2492)	<=	VN_out_sigd(691);
CN_in_sigd(2916)	<=	VN_out_sigd(691);
CN_in_sigd(4332)	<=	VN_out_sigd(691);
CN_in_sigd(1252)	<=	VN_out_sigd(692);
CN_in_sigd(2500)	<=	VN_out_sigd(692);
CN_in_sigd(2924)	<=	VN_out_sigd(692);
CN_in_sigd(4340)	<=	VN_out_sigd(692);
CN_in_sigd(1260)	<=	VN_out_sigd(693);
CN_in_sigd(2508)	<=	VN_out_sigd(693);
CN_in_sigd(2932)	<=	VN_out_sigd(693);
CN_in_sigd(4348)	<=	VN_out_sigd(693);
CN_in_sigd(1268)	<=	VN_out_sigd(694);
CN_in_sigd(2516)	<=	VN_out_sigd(694);
CN_in_sigd(2940)	<=	VN_out_sigd(694);
CN_in_sigd(4356)	<=	VN_out_sigd(694);
CN_in_sigd(1276)	<=	VN_out_sigd(695);
CN_in_sigd(2524)	<=	VN_out_sigd(695);
CN_in_sigd(2948)	<=	VN_out_sigd(695);
CN_in_sigd(4364)	<=	VN_out_sigd(695);
CN_in_sigd(1284)	<=	VN_out_sigd(696);
CN_in_sigd(2532)	<=	VN_out_sigd(696);
CN_in_sigd(2956)	<=	VN_out_sigd(696);
CN_in_sigd(4372)	<=	VN_out_sigd(696);
CN_in_sigd(1292)	<=	VN_out_sigd(697);
CN_in_sigd(2540)	<=	VN_out_sigd(697);
CN_in_sigd(2964)	<=	VN_out_sigd(697);
CN_in_sigd(4380)	<=	VN_out_sigd(697);
CN_in_sigd(868)	<=	VN_out_sigd(698);
CN_in_sigd(2548)	<=	VN_out_sigd(698);
CN_in_sigd(2972)	<=	VN_out_sigd(698);
CN_in_sigd(4388)	<=	VN_out_sigd(698);
CN_in_sigd(876)	<=	VN_out_sigd(699);
CN_in_sigd(2556)	<=	VN_out_sigd(699);
CN_in_sigd(2980)	<=	VN_out_sigd(699);
CN_in_sigd(4396)	<=	VN_out_sigd(699);
CN_in_sigd(884)	<=	VN_out_sigd(700);
CN_in_sigd(2564)	<=	VN_out_sigd(700);
CN_in_sigd(2988)	<=	VN_out_sigd(700);
CN_in_sigd(4404)	<=	VN_out_sigd(700);
CN_in_sigd(892)	<=	VN_out_sigd(701);
CN_in_sigd(2572)	<=	VN_out_sigd(701);
CN_in_sigd(2996)	<=	VN_out_sigd(701);
CN_in_sigd(4412)	<=	VN_out_sigd(701);
CN_in_sigd(84)	<=	VN_out_sigd(702);
CN_in_sigd(1628)	<=	VN_out_sigd(702);
CN_in_sigd(3740)	<=	VN_out_sigd(702);
CN_in_sigd(4820)	<=	VN_out_sigd(702);
CN_in_sigd(92)	<=	VN_out_sigd(703);
CN_in_sigd(1636)	<=	VN_out_sigd(703);
CN_in_sigd(3748)	<=	VN_out_sigd(703);
CN_in_sigd(4828)	<=	VN_out_sigd(703);
CN_in_sigd(100)	<=	VN_out_sigd(704);
CN_in_sigd(1644)	<=	VN_out_sigd(704);
CN_in_sigd(3756)	<=	VN_out_sigd(704);
CN_in_sigd(4836)	<=	VN_out_sigd(704);
CN_in_sigd(108)	<=	VN_out_sigd(705);
CN_in_sigd(1652)	<=	VN_out_sigd(705);
CN_in_sigd(3764)	<=	VN_out_sigd(705);
CN_in_sigd(4844)	<=	VN_out_sigd(705);
CN_in_sigd(116)	<=	VN_out_sigd(706);
CN_in_sigd(1660)	<=	VN_out_sigd(706);
CN_in_sigd(3772)	<=	VN_out_sigd(706);
CN_in_sigd(4852)	<=	VN_out_sigd(706);
CN_in_sigd(124)	<=	VN_out_sigd(707);
CN_in_sigd(1668)	<=	VN_out_sigd(707);
CN_in_sigd(3780)	<=	VN_out_sigd(707);
CN_in_sigd(4860)	<=	VN_out_sigd(707);
CN_in_sigd(132)	<=	VN_out_sigd(708);
CN_in_sigd(1676)	<=	VN_out_sigd(708);
CN_in_sigd(3788)	<=	VN_out_sigd(708);
CN_in_sigd(4868)	<=	VN_out_sigd(708);
CN_in_sigd(140)	<=	VN_out_sigd(709);
CN_in_sigd(1684)	<=	VN_out_sigd(709);
CN_in_sigd(3796)	<=	VN_out_sigd(709);
CN_in_sigd(4876)	<=	VN_out_sigd(709);
CN_in_sigd(148)	<=	VN_out_sigd(710);
CN_in_sigd(1692)	<=	VN_out_sigd(710);
CN_in_sigd(3804)	<=	VN_out_sigd(710);
CN_in_sigd(4884)	<=	VN_out_sigd(710);
CN_in_sigd(156)	<=	VN_out_sigd(711);
CN_in_sigd(1700)	<=	VN_out_sigd(711);
CN_in_sigd(3812)	<=	VN_out_sigd(711);
CN_in_sigd(4892)	<=	VN_out_sigd(711);
CN_in_sigd(164)	<=	VN_out_sigd(712);
CN_in_sigd(1708)	<=	VN_out_sigd(712);
CN_in_sigd(3820)	<=	VN_out_sigd(712);
CN_in_sigd(4900)	<=	VN_out_sigd(712);
CN_in_sigd(172)	<=	VN_out_sigd(713);
CN_in_sigd(1716)	<=	VN_out_sigd(713);
CN_in_sigd(3828)	<=	VN_out_sigd(713);
CN_in_sigd(4908)	<=	VN_out_sigd(713);
CN_in_sigd(180)	<=	VN_out_sigd(714);
CN_in_sigd(1724)	<=	VN_out_sigd(714);
CN_in_sigd(3836)	<=	VN_out_sigd(714);
CN_in_sigd(4916)	<=	VN_out_sigd(714);
CN_in_sigd(188)	<=	VN_out_sigd(715);
CN_in_sigd(1300)	<=	VN_out_sigd(715);
CN_in_sigd(3844)	<=	VN_out_sigd(715);
CN_in_sigd(4924)	<=	VN_out_sigd(715);
CN_in_sigd(196)	<=	VN_out_sigd(716);
CN_in_sigd(1308)	<=	VN_out_sigd(716);
CN_in_sigd(3852)	<=	VN_out_sigd(716);
CN_in_sigd(4932)	<=	VN_out_sigd(716);
CN_in_sigd(204)	<=	VN_out_sigd(717);
CN_in_sigd(1316)	<=	VN_out_sigd(717);
CN_in_sigd(3860)	<=	VN_out_sigd(717);
CN_in_sigd(4940)	<=	VN_out_sigd(717);
CN_in_sigd(212)	<=	VN_out_sigd(718);
CN_in_sigd(1324)	<=	VN_out_sigd(718);
CN_in_sigd(3868)	<=	VN_out_sigd(718);
CN_in_sigd(4948)	<=	VN_out_sigd(718);
CN_in_sigd(220)	<=	VN_out_sigd(719);
CN_in_sigd(1332)	<=	VN_out_sigd(719);
CN_in_sigd(3876)	<=	VN_out_sigd(719);
CN_in_sigd(4956)	<=	VN_out_sigd(719);
CN_in_sigd(228)	<=	VN_out_sigd(720);
CN_in_sigd(1340)	<=	VN_out_sigd(720);
CN_in_sigd(3884)	<=	VN_out_sigd(720);
CN_in_sigd(4964)	<=	VN_out_sigd(720);
CN_in_sigd(236)	<=	VN_out_sigd(721);
CN_in_sigd(1348)	<=	VN_out_sigd(721);
CN_in_sigd(3460)	<=	VN_out_sigd(721);
CN_in_sigd(4972)	<=	VN_out_sigd(721);
CN_in_sigd(244)	<=	VN_out_sigd(722);
CN_in_sigd(1356)	<=	VN_out_sigd(722);
CN_in_sigd(3468)	<=	VN_out_sigd(722);
CN_in_sigd(4980)	<=	VN_out_sigd(722);
CN_in_sigd(252)	<=	VN_out_sigd(723);
CN_in_sigd(1364)	<=	VN_out_sigd(723);
CN_in_sigd(3476)	<=	VN_out_sigd(723);
CN_in_sigd(4988)	<=	VN_out_sigd(723);
CN_in_sigd(260)	<=	VN_out_sigd(724);
CN_in_sigd(1372)	<=	VN_out_sigd(724);
CN_in_sigd(3484)	<=	VN_out_sigd(724);
CN_in_sigd(4996)	<=	VN_out_sigd(724);
CN_in_sigd(268)	<=	VN_out_sigd(725);
CN_in_sigd(1380)	<=	VN_out_sigd(725);
CN_in_sigd(3492)	<=	VN_out_sigd(725);
CN_in_sigd(5004)	<=	VN_out_sigd(725);
CN_in_sigd(276)	<=	VN_out_sigd(726);
CN_in_sigd(1388)	<=	VN_out_sigd(726);
CN_in_sigd(3500)	<=	VN_out_sigd(726);
CN_in_sigd(5012)	<=	VN_out_sigd(726);
CN_in_sigd(284)	<=	VN_out_sigd(727);
CN_in_sigd(1396)	<=	VN_out_sigd(727);
CN_in_sigd(3508)	<=	VN_out_sigd(727);
CN_in_sigd(5020)	<=	VN_out_sigd(727);
CN_in_sigd(292)	<=	VN_out_sigd(728);
CN_in_sigd(1404)	<=	VN_out_sigd(728);
CN_in_sigd(3516)	<=	VN_out_sigd(728);
CN_in_sigd(5028)	<=	VN_out_sigd(728);
CN_in_sigd(300)	<=	VN_out_sigd(729);
CN_in_sigd(1412)	<=	VN_out_sigd(729);
CN_in_sigd(3524)	<=	VN_out_sigd(729);
CN_in_sigd(5036)	<=	VN_out_sigd(729);
CN_in_sigd(308)	<=	VN_out_sigd(730);
CN_in_sigd(1420)	<=	VN_out_sigd(730);
CN_in_sigd(3532)	<=	VN_out_sigd(730);
CN_in_sigd(5044)	<=	VN_out_sigd(730);
CN_in_sigd(316)	<=	VN_out_sigd(731);
CN_in_sigd(1428)	<=	VN_out_sigd(731);
CN_in_sigd(3540)	<=	VN_out_sigd(731);
CN_in_sigd(5052)	<=	VN_out_sigd(731);
CN_in_sigd(324)	<=	VN_out_sigd(732);
CN_in_sigd(1436)	<=	VN_out_sigd(732);
CN_in_sigd(3548)	<=	VN_out_sigd(732);
CN_in_sigd(5060)	<=	VN_out_sigd(732);
CN_in_sigd(332)	<=	VN_out_sigd(733);
CN_in_sigd(1444)	<=	VN_out_sigd(733);
CN_in_sigd(3556)	<=	VN_out_sigd(733);
CN_in_sigd(5068)	<=	VN_out_sigd(733);
CN_in_sigd(340)	<=	VN_out_sigd(734);
CN_in_sigd(1452)	<=	VN_out_sigd(734);
CN_in_sigd(3564)	<=	VN_out_sigd(734);
CN_in_sigd(5076)	<=	VN_out_sigd(734);
CN_in_sigd(348)	<=	VN_out_sigd(735);
CN_in_sigd(1460)	<=	VN_out_sigd(735);
CN_in_sigd(3572)	<=	VN_out_sigd(735);
CN_in_sigd(5084)	<=	VN_out_sigd(735);
CN_in_sigd(356)	<=	VN_out_sigd(736);
CN_in_sigd(1468)	<=	VN_out_sigd(736);
CN_in_sigd(3580)	<=	VN_out_sigd(736);
CN_in_sigd(5092)	<=	VN_out_sigd(736);
CN_in_sigd(364)	<=	VN_out_sigd(737);
CN_in_sigd(1476)	<=	VN_out_sigd(737);
CN_in_sigd(3588)	<=	VN_out_sigd(737);
CN_in_sigd(5100)	<=	VN_out_sigd(737);
CN_in_sigd(372)	<=	VN_out_sigd(738);
CN_in_sigd(1484)	<=	VN_out_sigd(738);
CN_in_sigd(3596)	<=	VN_out_sigd(738);
CN_in_sigd(5108)	<=	VN_out_sigd(738);
CN_in_sigd(380)	<=	VN_out_sigd(739);
CN_in_sigd(1492)	<=	VN_out_sigd(739);
CN_in_sigd(3604)	<=	VN_out_sigd(739);
CN_in_sigd(5116)	<=	VN_out_sigd(739);
CN_in_sigd(388)	<=	VN_out_sigd(740);
CN_in_sigd(1500)	<=	VN_out_sigd(740);
CN_in_sigd(3612)	<=	VN_out_sigd(740);
CN_in_sigd(5124)	<=	VN_out_sigd(740);
CN_in_sigd(396)	<=	VN_out_sigd(741);
CN_in_sigd(1508)	<=	VN_out_sigd(741);
CN_in_sigd(3620)	<=	VN_out_sigd(741);
CN_in_sigd(5132)	<=	VN_out_sigd(741);
CN_in_sigd(404)	<=	VN_out_sigd(742);
CN_in_sigd(1516)	<=	VN_out_sigd(742);
CN_in_sigd(3628)	<=	VN_out_sigd(742);
CN_in_sigd(5140)	<=	VN_out_sigd(742);
CN_in_sigd(412)	<=	VN_out_sigd(743);
CN_in_sigd(1524)	<=	VN_out_sigd(743);
CN_in_sigd(3636)	<=	VN_out_sigd(743);
CN_in_sigd(5148)	<=	VN_out_sigd(743);
CN_in_sigd(420)	<=	VN_out_sigd(744);
CN_in_sigd(1532)	<=	VN_out_sigd(744);
CN_in_sigd(3644)	<=	VN_out_sigd(744);
CN_in_sigd(5156)	<=	VN_out_sigd(744);
CN_in_sigd(428)	<=	VN_out_sigd(745);
CN_in_sigd(1540)	<=	VN_out_sigd(745);
CN_in_sigd(3652)	<=	VN_out_sigd(745);
CN_in_sigd(5164)	<=	VN_out_sigd(745);
CN_in_sigd(4)	<=	VN_out_sigd(746);
CN_in_sigd(1548)	<=	VN_out_sigd(746);
CN_in_sigd(3660)	<=	VN_out_sigd(746);
CN_in_sigd(5172)	<=	VN_out_sigd(746);
CN_in_sigd(12)	<=	VN_out_sigd(747);
CN_in_sigd(1556)	<=	VN_out_sigd(747);
CN_in_sigd(3668)	<=	VN_out_sigd(747);
CN_in_sigd(5180)	<=	VN_out_sigd(747);
CN_in_sigd(20)	<=	VN_out_sigd(748);
CN_in_sigd(1564)	<=	VN_out_sigd(748);
CN_in_sigd(3676)	<=	VN_out_sigd(748);
CN_in_sigd(4756)	<=	VN_out_sigd(748);
CN_in_sigd(28)	<=	VN_out_sigd(749);
CN_in_sigd(1572)	<=	VN_out_sigd(749);
CN_in_sigd(3684)	<=	VN_out_sigd(749);
CN_in_sigd(4764)	<=	VN_out_sigd(749);
CN_in_sigd(36)	<=	VN_out_sigd(750);
CN_in_sigd(1580)	<=	VN_out_sigd(750);
CN_in_sigd(3692)	<=	VN_out_sigd(750);
CN_in_sigd(4772)	<=	VN_out_sigd(750);
CN_in_sigd(44)	<=	VN_out_sigd(751);
CN_in_sigd(1588)	<=	VN_out_sigd(751);
CN_in_sigd(3700)	<=	VN_out_sigd(751);
CN_in_sigd(4780)	<=	VN_out_sigd(751);
CN_in_sigd(52)	<=	VN_out_sigd(752);
CN_in_sigd(1596)	<=	VN_out_sigd(752);
CN_in_sigd(3708)	<=	VN_out_sigd(752);
CN_in_sigd(4788)	<=	VN_out_sigd(752);
CN_in_sigd(60)	<=	VN_out_sigd(753);
CN_in_sigd(1604)	<=	VN_out_sigd(753);
CN_in_sigd(3716)	<=	VN_out_sigd(753);
CN_in_sigd(4796)	<=	VN_out_sigd(753);
CN_in_sigd(68)	<=	VN_out_sigd(754);
CN_in_sigd(1612)	<=	VN_out_sigd(754);
CN_in_sigd(3724)	<=	VN_out_sigd(754);
CN_in_sigd(4804)	<=	VN_out_sigd(754);
CN_in_sigd(76)	<=	VN_out_sigd(755);
CN_in_sigd(1620)	<=	VN_out_sigd(755);
CN_in_sigd(3732)	<=	VN_out_sigd(755);
CN_in_sigd(4812)	<=	VN_out_sigd(755);
CN_in_sigd(580)	<=	VN_out_sigd(756);
CN_in_sigd(2132)	<=	VN_out_sigd(756);
CN_in_sigd(3084)	<=	VN_out_sigd(756);
CN_in_sigd(4084)	<=	VN_out_sigd(756);
CN_in_sigd(588)	<=	VN_out_sigd(757);
CN_in_sigd(2140)	<=	VN_out_sigd(757);
CN_in_sigd(3092)	<=	VN_out_sigd(757);
CN_in_sigd(4092)	<=	VN_out_sigd(757);
CN_in_sigd(596)	<=	VN_out_sigd(758);
CN_in_sigd(2148)	<=	VN_out_sigd(758);
CN_in_sigd(3100)	<=	VN_out_sigd(758);
CN_in_sigd(4100)	<=	VN_out_sigd(758);
CN_in_sigd(604)	<=	VN_out_sigd(759);
CN_in_sigd(2156)	<=	VN_out_sigd(759);
CN_in_sigd(3108)	<=	VN_out_sigd(759);
CN_in_sigd(4108)	<=	VN_out_sigd(759);
CN_in_sigd(612)	<=	VN_out_sigd(760);
CN_in_sigd(1732)	<=	VN_out_sigd(760);
CN_in_sigd(3116)	<=	VN_out_sigd(760);
CN_in_sigd(4116)	<=	VN_out_sigd(760);
CN_in_sigd(620)	<=	VN_out_sigd(761);
CN_in_sigd(1740)	<=	VN_out_sigd(761);
CN_in_sigd(3124)	<=	VN_out_sigd(761);
CN_in_sigd(4124)	<=	VN_out_sigd(761);
CN_in_sigd(628)	<=	VN_out_sigd(762);
CN_in_sigd(1748)	<=	VN_out_sigd(762);
CN_in_sigd(3132)	<=	VN_out_sigd(762);
CN_in_sigd(4132)	<=	VN_out_sigd(762);
CN_in_sigd(636)	<=	VN_out_sigd(763);
CN_in_sigd(1756)	<=	VN_out_sigd(763);
CN_in_sigd(3140)	<=	VN_out_sigd(763);
CN_in_sigd(4140)	<=	VN_out_sigd(763);
CN_in_sigd(644)	<=	VN_out_sigd(764);
CN_in_sigd(1764)	<=	VN_out_sigd(764);
CN_in_sigd(3148)	<=	VN_out_sigd(764);
CN_in_sigd(4148)	<=	VN_out_sigd(764);
CN_in_sigd(652)	<=	VN_out_sigd(765);
CN_in_sigd(1772)	<=	VN_out_sigd(765);
CN_in_sigd(3156)	<=	VN_out_sigd(765);
CN_in_sigd(4156)	<=	VN_out_sigd(765);
CN_in_sigd(660)	<=	VN_out_sigd(766);
CN_in_sigd(1780)	<=	VN_out_sigd(766);
CN_in_sigd(3164)	<=	VN_out_sigd(766);
CN_in_sigd(4164)	<=	VN_out_sigd(766);
CN_in_sigd(668)	<=	VN_out_sigd(767);
CN_in_sigd(1788)	<=	VN_out_sigd(767);
CN_in_sigd(3172)	<=	VN_out_sigd(767);
CN_in_sigd(4172)	<=	VN_out_sigd(767);
CN_in_sigd(676)	<=	VN_out_sigd(768);
CN_in_sigd(1796)	<=	VN_out_sigd(768);
CN_in_sigd(3180)	<=	VN_out_sigd(768);
CN_in_sigd(4180)	<=	VN_out_sigd(768);
CN_in_sigd(684)	<=	VN_out_sigd(769);
CN_in_sigd(1804)	<=	VN_out_sigd(769);
CN_in_sigd(3188)	<=	VN_out_sigd(769);
CN_in_sigd(4188)	<=	VN_out_sigd(769);
CN_in_sigd(692)	<=	VN_out_sigd(770);
CN_in_sigd(1812)	<=	VN_out_sigd(770);
CN_in_sigd(3196)	<=	VN_out_sigd(770);
CN_in_sigd(4196)	<=	VN_out_sigd(770);
CN_in_sigd(700)	<=	VN_out_sigd(771);
CN_in_sigd(1820)	<=	VN_out_sigd(771);
CN_in_sigd(3204)	<=	VN_out_sigd(771);
CN_in_sigd(4204)	<=	VN_out_sigd(771);
CN_in_sigd(708)	<=	VN_out_sigd(772);
CN_in_sigd(1828)	<=	VN_out_sigd(772);
CN_in_sigd(3212)	<=	VN_out_sigd(772);
CN_in_sigd(4212)	<=	VN_out_sigd(772);
CN_in_sigd(716)	<=	VN_out_sigd(773);
CN_in_sigd(1836)	<=	VN_out_sigd(773);
CN_in_sigd(3220)	<=	VN_out_sigd(773);
CN_in_sigd(4220)	<=	VN_out_sigd(773);
CN_in_sigd(724)	<=	VN_out_sigd(774);
CN_in_sigd(1844)	<=	VN_out_sigd(774);
CN_in_sigd(3228)	<=	VN_out_sigd(774);
CN_in_sigd(4228)	<=	VN_out_sigd(774);
CN_in_sigd(732)	<=	VN_out_sigd(775);
CN_in_sigd(1852)	<=	VN_out_sigd(775);
CN_in_sigd(3236)	<=	VN_out_sigd(775);
CN_in_sigd(4236)	<=	VN_out_sigd(775);
CN_in_sigd(740)	<=	VN_out_sigd(776);
CN_in_sigd(1860)	<=	VN_out_sigd(776);
CN_in_sigd(3244)	<=	VN_out_sigd(776);
CN_in_sigd(4244)	<=	VN_out_sigd(776);
CN_in_sigd(748)	<=	VN_out_sigd(777);
CN_in_sigd(1868)	<=	VN_out_sigd(777);
CN_in_sigd(3252)	<=	VN_out_sigd(777);
CN_in_sigd(4252)	<=	VN_out_sigd(777);
CN_in_sigd(756)	<=	VN_out_sigd(778);
CN_in_sigd(1876)	<=	VN_out_sigd(778);
CN_in_sigd(3260)	<=	VN_out_sigd(778);
CN_in_sigd(4260)	<=	VN_out_sigd(778);
CN_in_sigd(764)	<=	VN_out_sigd(779);
CN_in_sigd(1884)	<=	VN_out_sigd(779);
CN_in_sigd(3268)	<=	VN_out_sigd(779);
CN_in_sigd(4268)	<=	VN_out_sigd(779);
CN_in_sigd(772)	<=	VN_out_sigd(780);
CN_in_sigd(1892)	<=	VN_out_sigd(780);
CN_in_sigd(3276)	<=	VN_out_sigd(780);
CN_in_sigd(4276)	<=	VN_out_sigd(780);
CN_in_sigd(780)	<=	VN_out_sigd(781);
CN_in_sigd(1900)	<=	VN_out_sigd(781);
CN_in_sigd(3284)	<=	VN_out_sigd(781);
CN_in_sigd(4284)	<=	VN_out_sigd(781);
CN_in_sigd(788)	<=	VN_out_sigd(782);
CN_in_sigd(1908)	<=	VN_out_sigd(782);
CN_in_sigd(3292)	<=	VN_out_sigd(782);
CN_in_sigd(4292)	<=	VN_out_sigd(782);
CN_in_sigd(796)	<=	VN_out_sigd(783);
CN_in_sigd(1916)	<=	VN_out_sigd(783);
CN_in_sigd(3300)	<=	VN_out_sigd(783);
CN_in_sigd(4300)	<=	VN_out_sigd(783);
CN_in_sigd(804)	<=	VN_out_sigd(784);
CN_in_sigd(1924)	<=	VN_out_sigd(784);
CN_in_sigd(3308)	<=	VN_out_sigd(784);
CN_in_sigd(4308)	<=	VN_out_sigd(784);
CN_in_sigd(812)	<=	VN_out_sigd(785);
CN_in_sigd(1932)	<=	VN_out_sigd(785);
CN_in_sigd(3316)	<=	VN_out_sigd(785);
CN_in_sigd(4316)	<=	VN_out_sigd(785);
CN_in_sigd(820)	<=	VN_out_sigd(786);
CN_in_sigd(1940)	<=	VN_out_sigd(786);
CN_in_sigd(3324)	<=	VN_out_sigd(786);
CN_in_sigd(3892)	<=	VN_out_sigd(786);
CN_in_sigd(828)	<=	VN_out_sigd(787);
CN_in_sigd(1948)	<=	VN_out_sigd(787);
CN_in_sigd(3332)	<=	VN_out_sigd(787);
CN_in_sigd(3900)	<=	VN_out_sigd(787);
CN_in_sigd(836)	<=	VN_out_sigd(788);
CN_in_sigd(1956)	<=	VN_out_sigd(788);
CN_in_sigd(3340)	<=	VN_out_sigd(788);
CN_in_sigd(3908)	<=	VN_out_sigd(788);
CN_in_sigd(844)	<=	VN_out_sigd(789);
CN_in_sigd(1964)	<=	VN_out_sigd(789);
CN_in_sigd(3348)	<=	VN_out_sigd(789);
CN_in_sigd(3916)	<=	VN_out_sigd(789);
CN_in_sigd(852)	<=	VN_out_sigd(790);
CN_in_sigd(1972)	<=	VN_out_sigd(790);
CN_in_sigd(3356)	<=	VN_out_sigd(790);
CN_in_sigd(3924)	<=	VN_out_sigd(790);
CN_in_sigd(860)	<=	VN_out_sigd(791);
CN_in_sigd(1980)	<=	VN_out_sigd(791);
CN_in_sigd(3364)	<=	VN_out_sigd(791);
CN_in_sigd(3932)	<=	VN_out_sigd(791);
CN_in_sigd(436)	<=	VN_out_sigd(792);
CN_in_sigd(1988)	<=	VN_out_sigd(792);
CN_in_sigd(3372)	<=	VN_out_sigd(792);
CN_in_sigd(3940)	<=	VN_out_sigd(792);
CN_in_sigd(444)	<=	VN_out_sigd(793);
CN_in_sigd(1996)	<=	VN_out_sigd(793);
CN_in_sigd(3380)	<=	VN_out_sigd(793);
CN_in_sigd(3948)	<=	VN_out_sigd(793);
CN_in_sigd(452)	<=	VN_out_sigd(794);
CN_in_sigd(2004)	<=	VN_out_sigd(794);
CN_in_sigd(3388)	<=	VN_out_sigd(794);
CN_in_sigd(3956)	<=	VN_out_sigd(794);
CN_in_sigd(460)	<=	VN_out_sigd(795);
CN_in_sigd(2012)	<=	VN_out_sigd(795);
CN_in_sigd(3396)	<=	VN_out_sigd(795);
CN_in_sigd(3964)	<=	VN_out_sigd(795);
CN_in_sigd(468)	<=	VN_out_sigd(796);
CN_in_sigd(2020)	<=	VN_out_sigd(796);
CN_in_sigd(3404)	<=	VN_out_sigd(796);
CN_in_sigd(3972)	<=	VN_out_sigd(796);
CN_in_sigd(476)	<=	VN_out_sigd(797);
CN_in_sigd(2028)	<=	VN_out_sigd(797);
CN_in_sigd(3412)	<=	VN_out_sigd(797);
CN_in_sigd(3980)	<=	VN_out_sigd(797);
CN_in_sigd(484)	<=	VN_out_sigd(798);
CN_in_sigd(2036)	<=	VN_out_sigd(798);
CN_in_sigd(3420)	<=	VN_out_sigd(798);
CN_in_sigd(3988)	<=	VN_out_sigd(798);
CN_in_sigd(492)	<=	VN_out_sigd(799);
CN_in_sigd(2044)	<=	VN_out_sigd(799);
CN_in_sigd(3428)	<=	VN_out_sigd(799);
CN_in_sigd(3996)	<=	VN_out_sigd(799);
CN_in_sigd(500)	<=	VN_out_sigd(800);
CN_in_sigd(2052)	<=	VN_out_sigd(800);
CN_in_sigd(3436)	<=	VN_out_sigd(800);
CN_in_sigd(4004)	<=	VN_out_sigd(800);
CN_in_sigd(508)	<=	VN_out_sigd(801);
CN_in_sigd(2060)	<=	VN_out_sigd(801);
CN_in_sigd(3444)	<=	VN_out_sigd(801);
CN_in_sigd(4012)	<=	VN_out_sigd(801);
CN_in_sigd(516)	<=	VN_out_sigd(802);
CN_in_sigd(2068)	<=	VN_out_sigd(802);
CN_in_sigd(3452)	<=	VN_out_sigd(802);
CN_in_sigd(4020)	<=	VN_out_sigd(802);
CN_in_sigd(524)	<=	VN_out_sigd(803);
CN_in_sigd(2076)	<=	VN_out_sigd(803);
CN_in_sigd(3028)	<=	VN_out_sigd(803);
CN_in_sigd(4028)	<=	VN_out_sigd(803);
CN_in_sigd(532)	<=	VN_out_sigd(804);
CN_in_sigd(2084)	<=	VN_out_sigd(804);
CN_in_sigd(3036)	<=	VN_out_sigd(804);
CN_in_sigd(4036)	<=	VN_out_sigd(804);
CN_in_sigd(540)	<=	VN_out_sigd(805);
CN_in_sigd(2092)	<=	VN_out_sigd(805);
CN_in_sigd(3044)	<=	VN_out_sigd(805);
CN_in_sigd(4044)	<=	VN_out_sigd(805);
CN_in_sigd(548)	<=	VN_out_sigd(806);
CN_in_sigd(2100)	<=	VN_out_sigd(806);
CN_in_sigd(3052)	<=	VN_out_sigd(806);
CN_in_sigd(4052)	<=	VN_out_sigd(806);
CN_in_sigd(556)	<=	VN_out_sigd(807);
CN_in_sigd(2108)	<=	VN_out_sigd(807);
CN_in_sigd(3060)	<=	VN_out_sigd(807);
CN_in_sigd(4060)	<=	VN_out_sigd(807);
CN_in_sigd(564)	<=	VN_out_sigd(808);
CN_in_sigd(2116)	<=	VN_out_sigd(808);
CN_in_sigd(3068)	<=	VN_out_sigd(808);
CN_in_sigd(4068)	<=	VN_out_sigd(808);
CN_in_sigd(572)	<=	VN_out_sigd(809);
CN_in_sigd(2124)	<=	VN_out_sigd(809);
CN_in_sigd(3076)	<=	VN_out_sigd(809);
CN_in_sigd(4076)	<=	VN_out_sigd(809);
CN_in_sigd(885)	<=	VN_out_sigd(810);
CN_in_sigd(2053)	<=	VN_out_sigd(810);
CN_in_sigd(2693)	<=	VN_out_sigd(810);
CN_in_sigd(4357)	<=	VN_out_sigd(810);
CN_in_sigd(893)	<=	VN_out_sigd(811);
CN_in_sigd(2061)	<=	VN_out_sigd(811);
CN_in_sigd(2701)	<=	VN_out_sigd(811);
CN_in_sigd(4365)	<=	VN_out_sigd(811);
CN_in_sigd(901)	<=	VN_out_sigd(812);
CN_in_sigd(2069)	<=	VN_out_sigd(812);
CN_in_sigd(2709)	<=	VN_out_sigd(812);
CN_in_sigd(4373)	<=	VN_out_sigd(812);
CN_in_sigd(909)	<=	VN_out_sigd(813);
CN_in_sigd(2077)	<=	VN_out_sigd(813);
CN_in_sigd(2717)	<=	VN_out_sigd(813);
CN_in_sigd(4381)	<=	VN_out_sigd(813);
CN_in_sigd(917)	<=	VN_out_sigd(814);
CN_in_sigd(2085)	<=	VN_out_sigd(814);
CN_in_sigd(2725)	<=	VN_out_sigd(814);
CN_in_sigd(4389)	<=	VN_out_sigd(814);
CN_in_sigd(925)	<=	VN_out_sigd(815);
CN_in_sigd(2093)	<=	VN_out_sigd(815);
CN_in_sigd(2733)	<=	VN_out_sigd(815);
CN_in_sigd(4397)	<=	VN_out_sigd(815);
CN_in_sigd(933)	<=	VN_out_sigd(816);
CN_in_sigd(2101)	<=	VN_out_sigd(816);
CN_in_sigd(2741)	<=	VN_out_sigd(816);
CN_in_sigd(4405)	<=	VN_out_sigd(816);
CN_in_sigd(941)	<=	VN_out_sigd(817);
CN_in_sigd(2109)	<=	VN_out_sigd(817);
CN_in_sigd(2749)	<=	VN_out_sigd(817);
CN_in_sigd(4413)	<=	VN_out_sigd(817);
CN_in_sigd(949)	<=	VN_out_sigd(818);
CN_in_sigd(2117)	<=	VN_out_sigd(818);
CN_in_sigd(2757)	<=	VN_out_sigd(818);
CN_in_sigd(4421)	<=	VN_out_sigd(818);
CN_in_sigd(957)	<=	VN_out_sigd(819);
CN_in_sigd(2125)	<=	VN_out_sigd(819);
CN_in_sigd(2765)	<=	VN_out_sigd(819);
CN_in_sigd(4429)	<=	VN_out_sigd(819);
CN_in_sigd(965)	<=	VN_out_sigd(820);
CN_in_sigd(2133)	<=	VN_out_sigd(820);
CN_in_sigd(2773)	<=	VN_out_sigd(820);
CN_in_sigd(4437)	<=	VN_out_sigd(820);
CN_in_sigd(973)	<=	VN_out_sigd(821);
CN_in_sigd(2141)	<=	VN_out_sigd(821);
CN_in_sigd(2781)	<=	VN_out_sigd(821);
CN_in_sigd(4445)	<=	VN_out_sigd(821);
CN_in_sigd(981)	<=	VN_out_sigd(822);
CN_in_sigd(2149)	<=	VN_out_sigd(822);
CN_in_sigd(2789)	<=	VN_out_sigd(822);
CN_in_sigd(4453)	<=	VN_out_sigd(822);
CN_in_sigd(989)	<=	VN_out_sigd(823);
CN_in_sigd(2157)	<=	VN_out_sigd(823);
CN_in_sigd(2797)	<=	VN_out_sigd(823);
CN_in_sigd(4461)	<=	VN_out_sigd(823);
CN_in_sigd(997)	<=	VN_out_sigd(824);
CN_in_sigd(1733)	<=	VN_out_sigd(824);
CN_in_sigd(2805)	<=	VN_out_sigd(824);
CN_in_sigd(4469)	<=	VN_out_sigd(824);
CN_in_sigd(1005)	<=	VN_out_sigd(825);
CN_in_sigd(1741)	<=	VN_out_sigd(825);
CN_in_sigd(2813)	<=	VN_out_sigd(825);
CN_in_sigd(4477)	<=	VN_out_sigd(825);
CN_in_sigd(1013)	<=	VN_out_sigd(826);
CN_in_sigd(1749)	<=	VN_out_sigd(826);
CN_in_sigd(2821)	<=	VN_out_sigd(826);
CN_in_sigd(4485)	<=	VN_out_sigd(826);
CN_in_sigd(1021)	<=	VN_out_sigd(827);
CN_in_sigd(1757)	<=	VN_out_sigd(827);
CN_in_sigd(2829)	<=	VN_out_sigd(827);
CN_in_sigd(4493)	<=	VN_out_sigd(827);
CN_in_sigd(1029)	<=	VN_out_sigd(828);
CN_in_sigd(1765)	<=	VN_out_sigd(828);
CN_in_sigd(2837)	<=	VN_out_sigd(828);
CN_in_sigd(4501)	<=	VN_out_sigd(828);
CN_in_sigd(1037)	<=	VN_out_sigd(829);
CN_in_sigd(1773)	<=	VN_out_sigd(829);
CN_in_sigd(2845)	<=	VN_out_sigd(829);
CN_in_sigd(4509)	<=	VN_out_sigd(829);
CN_in_sigd(1045)	<=	VN_out_sigd(830);
CN_in_sigd(1781)	<=	VN_out_sigd(830);
CN_in_sigd(2853)	<=	VN_out_sigd(830);
CN_in_sigd(4517)	<=	VN_out_sigd(830);
CN_in_sigd(1053)	<=	VN_out_sigd(831);
CN_in_sigd(1789)	<=	VN_out_sigd(831);
CN_in_sigd(2861)	<=	VN_out_sigd(831);
CN_in_sigd(4525)	<=	VN_out_sigd(831);
CN_in_sigd(1061)	<=	VN_out_sigd(832);
CN_in_sigd(1797)	<=	VN_out_sigd(832);
CN_in_sigd(2869)	<=	VN_out_sigd(832);
CN_in_sigd(4533)	<=	VN_out_sigd(832);
CN_in_sigd(1069)	<=	VN_out_sigd(833);
CN_in_sigd(1805)	<=	VN_out_sigd(833);
CN_in_sigd(2877)	<=	VN_out_sigd(833);
CN_in_sigd(4541)	<=	VN_out_sigd(833);
CN_in_sigd(1077)	<=	VN_out_sigd(834);
CN_in_sigd(1813)	<=	VN_out_sigd(834);
CN_in_sigd(2885)	<=	VN_out_sigd(834);
CN_in_sigd(4549)	<=	VN_out_sigd(834);
CN_in_sigd(1085)	<=	VN_out_sigd(835);
CN_in_sigd(1821)	<=	VN_out_sigd(835);
CN_in_sigd(2893)	<=	VN_out_sigd(835);
CN_in_sigd(4557)	<=	VN_out_sigd(835);
CN_in_sigd(1093)	<=	VN_out_sigd(836);
CN_in_sigd(1829)	<=	VN_out_sigd(836);
CN_in_sigd(2901)	<=	VN_out_sigd(836);
CN_in_sigd(4565)	<=	VN_out_sigd(836);
CN_in_sigd(1101)	<=	VN_out_sigd(837);
CN_in_sigd(1837)	<=	VN_out_sigd(837);
CN_in_sigd(2909)	<=	VN_out_sigd(837);
CN_in_sigd(4573)	<=	VN_out_sigd(837);
CN_in_sigd(1109)	<=	VN_out_sigd(838);
CN_in_sigd(1845)	<=	VN_out_sigd(838);
CN_in_sigd(2917)	<=	VN_out_sigd(838);
CN_in_sigd(4581)	<=	VN_out_sigd(838);
CN_in_sigd(1117)	<=	VN_out_sigd(839);
CN_in_sigd(1853)	<=	VN_out_sigd(839);
CN_in_sigd(2925)	<=	VN_out_sigd(839);
CN_in_sigd(4589)	<=	VN_out_sigd(839);
CN_in_sigd(1125)	<=	VN_out_sigd(840);
CN_in_sigd(1861)	<=	VN_out_sigd(840);
CN_in_sigd(2933)	<=	VN_out_sigd(840);
CN_in_sigd(4597)	<=	VN_out_sigd(840);
CN_in_sigd(1133)	<=	VN_out_sigd(841);
CN_in_sigd(1869)	<=	VN_out_sigd(841);
CN_in_sigd(2941)	<=	VN_out_sigd(841);
CN_in_sigd(4605)	<=	VN_out_sigd(841);
CN_in_sigd(1141)	<=	VN_out_sigd(842);
CN_in_sigd(1877)	<=	VN_out_sigd(842);
CN_in_sigd(2949)	<=	VN_out_sigd(842);
CN_in_sigd(4613)	<=	VN_out_sigd(842);
CN_in_sigd(1149)	<=	VN_out_sigd(843);
CN_in_sigd(1885)	<=	VN_out_sigd(843);
CN_in_sigd(2957)	<=	VN_out_sigd(843);
CN_in_sigd(4621)	<=	VN_out_sigd(843);
CN_in_sigd(1157)	<=	VN_out_sigd(844);
CN_in_sigd(1893)	<=	VN_out_sigd(844);
CN_in_sigd(2965)	<=	VN_out_sigd(844);
CN_in_sigd(4629)	<=	VN_out_sigd(844);
CN_in_sigd(1165)	<=	VN_out_sigd(845);
CN_in_sigd(1901)	<=	VN_out_sigd(845);
CN_in_sigd(2973)	<=	VN_out_sigd(845);
CN_in_sigd(4637)	<=	VN_out_sigd(845);
CN_in_sigd(1173)	<=	VN_out_sigd(846);
CN_in_sigd(1909)	<=	VN_out_sigd(846);
CN_in_sigd(2981)	<=	VN_out_sigd(846);
CN_in_sigd(4645)	<=	VN_out_sigd(846);
CN_in_sigd(1181)	<=	VN_out_sigd(847);
CN_in_sigd(1917)	<=	VN_out_sigd(847);
CN_in_sigd(2989)	<=	VN_out_sigd(847);
CN_in_sigd(4653)	<=	VN_out_sigd(847);
CN_in_sigd(1189)	<=	VN_out_sigd(848);
CN_in_sigd(1925)	<=	VN_out_sigd(848);
CN_in_sigd(2997)	<=	VN_out_sigd(848);
CN_in_sigd(4661)	<=	VN_out_sigd(848);
CN_in_sigd(1197)	<=	VN_out_sigd(849);
CN_in_sigd(1933)	<=	VN_out_sigd(849);
CN_in_sigd(3005)	<=	VN_out_sigd(849);
CN_in_sigd(4669)	<=	VN_out_sigd(849);
CN_in_sigd(1205)	<=	VN_out_sigd(850);
CN_in_sigd(1941)	<=	VN_out_sigd(850);
CN_in_sigd(3013)	<=	VN_out_sigd(850);
CN_in_sigd(4677)	<=	VN_out_sigd(850);
CN_in_sigd(1213)	<=	VN_out_sigd(851);
CN_in_sigd(1949)	<=	VN_out_sigd(851);
CN_in_sigd(3021)	<=	VN_out_sigd(851);
CN_in_sigd(4685)	<=	VN_out_sigd(851);
CN_in_sigd(1221)	<=	VN_out_sigd(852);
CN_in_sigd(1957)	<=	VN_out_sigd(852);
CN_in_sigd(2597)	<=	VN_out_sigd(852);
CN_in_sigd(4693)	<=	VN_out_sigd(852);
CN_in_sigd(1229)	<=	VN_out_sigd(853);
CN_in_sigd(1965)	<=	VN_out_sigd(853);
CN_in_sigd(2605)	<=	VN_out_sigd(853);
CN_in_sigd(4701)	<=	VN_out_sigd(853);
CN_in_sigd(1237)	<=	VN_out_sigd(854);
CN_in_sigd(1973)	<=	VN_out_sigd(854);
CN_in_sigd(2613)	<=	VN_out_sigd(854);
CN_in_sigd(4709)	<=	VN_out_sigd(854);
CN_in_sigd(1245)	<=	VN_out_sigd(855);
CN_in_sigd(1981)	<=	VN_out_sigd(855);
CN_in_sigd(2621)	<=	VN_out_sigd(855);
CN_in_sigd(4717)	<=	VN_out_sigd(855);
CN_in_sigd(1253)	<=	VN_out_sigd(856);
CN_in_sigd(1989)	<=	VN_out_sigd(856);
CN_in_sigd(2629)	<=	VN_out_sigd(856);
CN_in_sigd(4725)	<=	VN_out_sigd(856);
CN_in_sigd(1261)	<=	VN_out_sigd(857);
CN_in_sigd(1997)	<=	VN_out_sigd(857);
CN_in_sigd(2637)	<=	VN_out_sigd(857);
CN_in_sigd(4733)	<=	VN_out_sigd(857);
CN_in_sigd(1269)	<=	VN_out_sigd(858);
CN_in_sigd(2005)	<=	VN_out_sigd(858);
CN_in_sigd(2645)	<=	VN_out_sigd(858);
CN_in_sigd(4741)	<=	VN_out_sigd(858);
CN_in_sigd(1277)	<=	VN_out_sigd(859);
CN_in_sigd(2013)	<=	VN_out_sigd(859);
CN_in_sigd(2653)	<=	VN_out_sigd(859);
CN_in_sigd(4749)	<=	VN_out_sigd(859);
CN_in_sigd(1285)	<=	VN_out_sigd(860);
CN_in_sigd(2021)	<=	VN_out_sigd(860);
CN_in_sigd(2661)	<=	VN_out_sigd(860);
CN_in_sigd(4325)	<=	VN_out_sigd(860);
CN_in_sigd(1293)	<=	VN_out_sigd(861);
CN_in_sigd(2029)	<=	VN_out_sigd(861);
CN_in_sigd(2669)	<=	VN_out_sigd(861);
CN_in_sigd(4333)	<=	VN_out_sigd(861);
CN_in_sigd(869)	<=	VN_out_sigd(862);
CN_in_sigd(2037)	<=	VN_out_sigd(862);
CN_in_sigd(2677)	<=	VN_out_sigd(862);
CN_in_sigd(4341)	<=	VN_out_sigd(862);
CN_in_sigd(877)	<=	VN_out_sigd(863);
CN_in_sigd(2045)	<=	VN_out_sigd(863);
CN_in_sigd(2685)	<=	VN_out_sigd(863);
CN_in_sigd(4349)	<=	VN_out_sigd(863);
CN_in_sigd(85)	<=	VN_out_sigd(864);
CN_in_sigd(1517)	<=	VN_out_sigd(864);
CN_in_sigd(3853)	<=	VN_out_sigd(864);
CN_in_sigd(5093)	<=	VN_out_sigd(864);
CN_in_sigd(93)	<=	VN_out_sigd(865);
CN_in_sigd(1525)	<=	VN_out_sigd(865);
CN_in_sigd(3861)	<=	VN_out_sigd(865);
CN_in_sigd(5101)	<=	VN_out_sigd(865);
CN_in_sigd(101)	<=	VN_out_sigd(866);
CN_in_sigd(1533)	<=	VN_out_sigd(866);
CN_in_sigd(3869)	<=	VN_out_sigd(866);
CN_in_sigd(5109)	<=	VN_out_sigd(866);
CN_in_sigd(109)	<=	VN_out_sigd(867);
CN_in_sigd(1541)	<=	VN_out_sigd(867);
CN_in_sigd(3877)	<=	VN_out_sigd(867);
CN_in_sigd(5117)	<=	VN_out_sigd(867);
CN_in_sigd(117)	<=	VN_out_sigd(868);
CN_in_sigd(1549)	<=	VN_out_sigd(868);
CN_in_sigd(3885)	<=	VN_out_sigd(868);
CN_in_sigd(5125)	<=	VN_out_sigd(868);
CN_in_sigd(125)	<=	VN_out_sigd(869);
CN_in_sigd(1557)	<=	VN_out_sigd(869);
CN_in_sigd(3461)	<=	VN_out_sigd(869);
CN_in_sigd(5133)	<=	VN_out_sigd(869);
CN_in_sigd(133)	<=	VN_out_sigd(870);
CN_in_sigd(1565)	<=	VN_out_sigd(870);
CN_in_sigd(3469)	<=	VN_out_sigd(870);
CN_in_sigd(5141)	<=	VN_out_sigd(870);
CN_in_sigd(141)	<=	VN_out_sigd(871);
CN_in_sigd(1573)	<=	VN_out_sigd(871);
CN_in_sigd(3477)	<=	VN_out_sigd(871);
CN_in_sigd(5149)	<=	VN_out_sigd(871);
CN_in_sigd(149)	<=	VN_out_sigd(872);
CN_in_sigd(1581)	<=	VN_out_sigd(872);
CN_in_sigd(3485)	<=	VN_out_sigd(872);
CN_in_sigd(5157)	<=	VN_out_sigd(872);
CN_in_sigd(157)	<=	VN_out_sigd(873);
CN_in_sigd(1589)	<=	VN_out_sigd(873);
CN_in_sigd(3493)	<=	VN_out_sigd(873);
CN_in_sigd(5165)	<=	VN_out_sigd(873);
CN_in_sigd(165)	<=	VN_out_sigd(874);
CN_in_sigd(1597)	<=	VN_out_sigd(874);
CN_in_sigd(3501)	<=	VN_out_sigd(874);
CN_in_sigd(5173)	<=	VN_out_sigd(874);
CN_in_sigd(173)	<=	VN_out_sigd(875);
CN_in_sigd(1605)	<=	VN_out_sigd(875);
CN_in_sigd(3509)	<=	VN_out_sigd(875);
CN_in_sigd(5181)	<=	VN_out_sigd(875);
CN_in_sigd(181)	<=	VN_out_sigd(876);
CN_in_sigd(1613)	<=	VN_out_sigd(876);
CN_in_sigd(3517)	<=	VN_out_sigd(876);
CN_in_sigd(4757)	<=	VN_out_sigd(876);
CN_in_sigd(189)	<=	VN_out_sigd(877);
CN_in_sigd(1621)	<=	VN_out_sigd(877);
CN_in_sigd(3525)	<=	VN_out_sigd(877);
CN_in_sigd(4765)	<=	VN_out_sigd(877);
CN_in_sigd(197)	<=	VN_out_sigd(878);
CN_in_sigd(1629)	<=	VN_out_sigd(878);
CN_in_sigd(3533)	<=	VN_out_sigd(878);
CN_in_sigd(4773)	<=	VN_out_sigd(878);
CN_in_sigd(205)	<=	VN_out_sigd(879);
CN_in_sigd(1637)	<=	VN_out_sigd(879);
CN_in_sigd(3541)	<=	VN_out_sigd(879);
CN_in_sigd(4781)	<=	VN_out_sigd(879);
CN_in_sigd(213)	<=	VN_out_sigd(880);
CN_in_sigd(1645)	<=	VN_out_sigd(880);
CN_in_sigd(3549)	<=	VN_out_sigd(880);
CN_in_sigd(4789)	<=	VN_out_sigd(880);
CN_in_sigd(221)	<=	VN_out_sigd(881);
CN_in_sigd(1653)	<=	VN_out_sigd(881);
CN_in_sigd(3557)	<=	VN_out_sigd(881);
CN_in_sigd(4797)	<=	VN_out_sigd(881);
CN_in_sigd(229)	<=	VN_out_sigd(882);
CN_in_sigd(1661)	<=	VN_out_sigd(882);
CN_in_sigd(3565)	<=	VN_out_sigd(882);
CN_in_sigd(4805)	<=	VN_out_sigd(882);
CN_in_sigd(237)	<=	VN_out_sigd(883);
CN_in_sigd(1669)	<=	VN_out_sigd(883);
CN_in_sigd(3573)	<=	VN_out_sigd(883);
CN_in_sigd(4813)	<=	VN_out_sigd(883);
CN_in_sigd(245)	<=	VN_out_sigd(884);
CN_in_sigd(1677)	<=	VN_out_sigd(884);
CN_in_sigd(3581)	<=	VN_out_sigd(884);
CN_in_sigd(4821)	<=	VN_out_sigd(884);
CN_in_sigd(253)	<=	VN_out_sigd(885);
CN_in_sigd(1685)	<=	VN_out_sigd(885);
CN_in_sigd(3589)	<=	VN_out_sigd(885);
CN_in_sigd(4829)	<=	VN_out_sigd(885);
CN_in_sigd(261)	<=	VN_out_sigd(886);
CN_in_sigd(1693)	<=	VN_out_sigd(886);
CN_in_sigd(3597)	<=	VN_out_sigd(886);
CN_in_sigd(4837)	<=	VN_out_sigd(886);
CN_in_sigd(269)	<=	VN_out_sigd(887);
CN_in_sigd(1701)	<=	VN_out_sigd(887);
CN_in_sigd(3605)	<=	VN_out_sigd(887);
CN_in_sigd(4845)	<=	VN_out_sigd(887);
CN_in_sigd(277)	<=	VN_out_sigd(888);
CN_in_sigd(1709)	<=	VN_out_sigd(888);
CN_in_sigd(3613)	<=	VN_out_sigd(888);
CN_in_sigd(4853)	<=	VN_out_sigd(888);
CN_in_sigd(285)	<=	VN_out_sigd(889);
CN_in_sigd(1717)	<=	VN_out_sigd(889);
CN_in_sigd(3621)	<=	VN_out_sigd(889);
CN_in_sigd(4861)	<=	VN_out_sigd(889);
CN_in_sigd(293)	<=	VN_out_sigd(890);
CN_in_sigd(1725)	<=	VN_out_sigd(890);
CN_in_sigd(3629)	<=	VN_out_sigd(890);
CN_in_sigd(4869)	<=	VN_out_sigd(890);
CN_in_sigd(301)	<=	VN_out_sigd(891);
CN_in_sigd(1301)	<=	VN_out_sigd(891);
CN_in_sigd(3637)	<=	VN_out_sigd(891);
CN_in_sigd(4877)	<=	VN_out_sigd(891);
CN_in_sigd(309)	<=	VN_out_sigd(892);
CN_in_sigd(1309)	<=	VN_out_sigd(892);
CN_in_sigd(3645)	<=	VN_out_sigd(892);
CN_in_sigd(4885)	<=	VN_out_sigd(892);
CN_in_sigd(317)	<=	VN_out_sigd(893);
CN_in_sigd(1317)	<=	VN_out_sigd(893);
CN_in_sigd(3653)	<=	VN_out_sigd(893);
CN_in_sigd(4893)	<=	VN_out_sigd(893);
CN_in_sigd(325)	<=	VN_out_sigd(894);
CN_in_sigd(1325)	<=	VN_out_sigd(894);
CN_in_sigd(3661)	<=	VN_out_sigd(894);
CN_in_sigd(4901)	<=	VN_out_sigd(894);
CN_in_sigd(333)	<=	VN_out_sigd(895);
CN_in_sigd(1333)	<=	VN_out_sigd(895);
CN_in_sigd(3669)	<=	VN_out_sigd(895);
CN_in_sigd(4909)	<=	VN_out_sigd(895);
CN_in_sigd(341)	<=	VN_out_sigd(896);
CN_in_sigd(1341)	<=	VN_out_sigd(896);
CN_in_sigd(3677)	<=	VN_out_sigd(896);
CN_in_sigd(4917)	<=	VN_out_sigd(896);
CN_in_sigd(349)	<=	VN_out_sigd(897);
CN_in_sigd(1349)	<=	VN_out_sigd(897);
CN_in_sigd(3685)	<=	VN_out_sigd(897);
CN_in_sigd(4925)	<=	VN_out_sigd(897);
CN_in_sigd(357)	<=	VN_out_sigd(898);
CN_in_sigd(1357)	<=	VN_out_sigd(898);
CN_in_sigd(3693)	<=	VN_out_sigd(898);
CN_in_sigd(4933)	<=	VN_out_sigd(898);
CN_in_sigd(365)	<=	VN_out_sigd(899);
CN_in_sigd(1365)	<=	VN_out_sigd(899);
CN_in_sigd(3701)	<=	VN_out_sigd(899);
CN_in_sigd(4941)	<=	VN_out_sigd(899);
CN_in_sigd(373)	<=	VN_out_sigd(900);
CN_in_sigd(1373)	<=	VN_out_sigd(900);
CN_in_sigd(3709)	<=	VN_out_sigd(900);
CN_in_sigd(4949)	<=	VN_out_sigd(900);
CN_in_sigd(381)	<=	VN_out_sigd(901);
CN_in_sigd(1381)	<=	VN_out_sigd(901);
CN_in_sigd(3717)	<=	VN_out_sigd(901);
CN_in_sigd(4957)	<=	VN_out_sigd(901);
CN_in_sigd(389)	<=	VN_out_sigd(902);
CN_in_sigd(1389)	<=	VN_out_sigd(902);
CN_in_sigd(3725)	<=	VN_out_sigd(902);
CN_in_sigd(4965)	<=	VN_out_sigd(902);
CN_in_sigd(397)	<=	VN_out_sigd(903);
CN_in_sigd(1397)	<=	VN_out_sigd(903);
CN_in_sigd(3733)	<=	VN_out_sigd(903);
CN_in_sigd(4973)	<=	VN_out_sigd(903);
CN_in_sigd(405)	<=	VN_out_sigd(904);
CN_in_sigd(1405)	<=	VN_out_sigd(904);
CN_in_sigd(3741)	<=	VN_out_sigd(904);
CN_in_sigd(4981)	<=	VN_out_sigd(904);
CN_in_sigd(413)	<=	VN_out_sigd(905);
CN_in_sigd(1413)	<=	VN_out_sigd(905);
CN_in_sigd(3749)	<=	VN_out_sigd(905);
CN_in_sigd(4989)	<=	VN_out_sigd(905);
CN_in_sigd(421)	<=	VN_out_sigd(906);
CN_in_sigd(1421)	<=	VN_out_sigd(906);
CN_in_sigd(3757)	<=	VN_out_sigd(906);
CN_in_sigd(4997)	<=	VN_out_sigd(906);
CN_in_sigd(429)	<=	VN_out_sigd(907);
CN_in_sigd(1429)	<=	VN_out_sigd(907);
CN_in_sigd(3765)	<=	VN_out_sigd(907);
CN_in_sigd(5005)	<=	VN_out_sigd(907);
CN_in_sigd(5)	<=	VN_out_sigd(908);
CN_in_sigd(1437)	<=	VN_out_sigd(908);
CN_in_sigd(3773)	<=	VN_out_sigd(908);
CN_in_sigd(5013)	<=	VN_out_sigd(908);
CN_in_sigd(13)	<=	VN_out_sigd(909);
CN_in_sigd(1445)	<=	VN_out_sigd(909);
CN_in_sigd(3781)	<=	VN_out_sigd(909);
CN_in_sigd(5021)	<=	VN_out_sigd(909);
CN_in_sigd(21)	<=	VN_out_sigd(910);
CN_in_sigd(1453)	<=	VN_out_sigd(910);
CN_in_sigd(3789)	<=	VN_out_sigd(910);
CN_in_sigd(5029)	<=	VN_out_sigd(910);
CN_in_sigd(29)	<=	VN_out_sigd(911);
CN_in_sigd(1461)	<=	VN_out_sigd(911);
CN_in_sigd(3797)	<=	VN_out_sigd(911);
CN_in_sigd(5037)	<=	VN_out_sigd(911);
CN_in_sigd(37)	<=	VN_out_sigd(912);
CN_in_sigd(1469)	<=	VN_out_sigd(912);
CN_in_sigd(3805)	<=	VN_out_sigd(912);
CN_in_sigd(5045)	<=	VN_out_sigd(912);
CN_in_sigd(45)	<=	VN_out_sigd(913);
CN_in_sigd(1477)	<=	VN_out_sigd(913);
CN_in_sigd(3813)	<=	VN_out_sigd(913);
CN_in_sigd(5053)	<=	VN_out_sigd(913);
CN_in_sigd(53)	<=	VN_out_sigd(914);
CN_in_sigd(1485)	<=	VN_out_sigd(914);
CN_in_sigd(3821)	<=	VN_out_sigd(914);
CN_in_sigd(5061)	<=	VN_out_sigd(914);
CN_in_sigd(61)	<=	VN_out_sigd(915);
CN_in_sigd(1493)	<=	VN_out_sigd(915);
CN_in_sigd(3829)	<=	VN_out_sigd(915);
CN_in_sigd(5069)	<=	VN_out_sigd(915);
CN_in_sigd(69)	<=	VN_out_sigd(916);
CN_in_sigd(1501)	<=	VN_out_sigd(916);
CN_in_sigd(3837)	<=	VN_out_sigd(916);
CN_in_sigd(5077)	<=	VN_out_sigd(916);
CN_in_sigd(77)	<=	VN_out_sigd(917);
CN_in_sigd(1509)	<=	VN_out_sigd(917);
CN_in_sigd(3845)	<=	VN_out_sigd(917);
CN_in_sigd(5085)	<=	VN_out_sigd(917);
CN_in_sigd(597)	<=	VN_out_sigd(918);
CN_in_sigd(2445)	<=	VN_out_sigd(918);
CN_in_sigd(3237)	<=	VN_out_sigd(918);
CN_in_sigd(4285)	<=	VN_out_sigd(918);
CN_in_sigd(605)	<=	VN_out_sigd(919);
CN_in_sigd(2453)	<=	VN_out_sigd(919);
CN_in_sigd(3245)	<=	VN_out_sigd(919);
CN_in_sigd(4293)	<=	VN_out_sigd(919);
CN_in_sigd(613)	<=	VN_out_sigd(920);
CN_in_sigd(2461)	<=	VN_out_sigd(920);
CN_in_sigd(3253)	<=	VN_out_sigd(920);
CN_in_sigd(4301)	<=	VN_out_sigd(920);
CN_in_sigd(621)	<=	VN_out_sigd(921);
CN_in_sigd(2469)	<=	VN_out_sigd(921);
CN_in_sigd(3261)	<=	VN_out_sigd(921);
CN_in_sigd(4309)	<=	VN_out_sigd(921);
CN_in_sigd(629)	<=	VN_out_sigd(922);
CN_in_sigd(2477)	<=	VN_out_sigd(922);
CN_in_sigd(3269)	<=	VN_out_sigd(922);
CN_in_sigd(4317)	<=	VN_out_sigd(922);
CN_in_sigd(637)	<=	VN_out_sigd(923);
CN_in_sigd(2485)	<=	VN_out_sigd(923);
CN_in_sigd(3277)	<=	VN_out_sigd(923);
CN_in_sigd(3893)	<=	VN_out_sigd(923);
CN_in_sigd(645)	<=	VN_out_sigd(924);
CN_in_sigd(2493)	<=	VN_out_sigd(924);
CN_in_sigd(3285)	<=	VN_out_sigd(924);
CN_in_sigd(3901)	<=	VN_out_sigd(924);
CN_in_sigd(653)	<=	VN_out_sigd(925);
CN_in_sigd(2501)	<=	VN_out_sigd(925);
CN_in_sigd(3293)	<=	VN_out_sigd(925);
CN_in_sigd(3909)	<=	VN_out_sigd(925);
CN_in_sigd(661)	<=	VN_out_sigd(926);
CN_in_sigd(2509)	<=	VN_out_sigd(926);
CN_in_sigd(3301)	<=	VN_out_sigd(926);
CN_in_sigd(3917)	<=	VN_out_sigd(926);
CN_in_sigd(669)	<=	VN_out_sigd(927);
CN_in_sigd(2517)	<=	VN_out_sigd(927);
CN_in_sigd(3309)	<=	VN_out_sigd(927);
CN_in_sigd(3925)	<=	VN_out_sigd(927);
CN_in_sigd(677)	<=	VN_out_sigd(928);
CN_in_sigd(2525)	<=	VN_out_sigd(928);
CN_in_sigd(3317)	<=	VN_out_sigd(928);
CN_in_sigd(3933)	<=	VN_out_sigd(928);
CN_in_sigd(685)	<=	VN_out_sigd(929);
CN_in_sigd(2533)	<=	VN_out_sigd(929);
CN_in_sigd(3325)	<=	VN_out_sigd(929);
CN_in_sigd(3941)	<=	VN_out_sigd(929);
CN_in_sigd(693)	<=	VN_out_sigd(930);
CN_in_sigd(2541)	<=	VN_out_sigd(930);
CN_in_sigd(3333)	<=	VN_out_sigd(930);
CN_in_sigd(3949)	<=	VN_out_sigd(930);
CN_in_sigd(701)	<=	VN_out_sigd(931);
CN_in_sigd(2549)	<=	VN_out_sigd(931);
CN_in_sigd(3341)	<=	VN_out_sigd(931);
CN_in_sigd(3957)	<=	VN_out_sigd(931);
CN_in_sigd(709)	<=	VN_out_sigd(932);
CN_in_sigd(2557)	<=	VN_out_sigd(932);
CN_in_sigd(3349)	<=	VN_out_sigd(932);
CN_in_sigd(3965)	<=	VN_out_sigd(932);
CN_in_sigd(717)	<=	VN_out_sigd(933);
CN_in_sigd(2565)	<=	VN_out_sigd(933);
CN_in_sigd(3357)	<=	VN_out_sigd(933);
CN_in_sigd(3973)	<=	VN_out_sigd(933);
CN_in_sigd(725)	<=	VN_out_sigd(934);
CN_in_sigd(2573)	<=	VN_out_sigd(934);
CN_in_sigd(3365)	<=	VN_out_sigd(934);
CN_in_sigd(3981)	<=	VN_out_sigd(934);
CN_in_sigd(733)	<=	VN_out_sigd(935);
CN_in_sigd(2581)	<=	VN_out_sigd(935);
CN_in_sigd(3373)	<=	VN_out_sigd(935);
CN_in_sigd(3989)	<=	VN_out_sigd(935);
CN_in_sigd(741)	<=	VN_out_sigd(936);
CN_in_sigd(2589)	<=	VN_out_sigd(936);
CN_in_sigd(3381)	<=	VN_out_sigd(936);
CN_in_sigd(3997)	<=	VN_out_sigd(936);
CN_in_sigd(749)	<=	VN_out_sigd(937);
CN_in_sigd(2165)	<=	VN_out_sigd(937);
CN_in_sigd(3389)	<=	VN_out_sigd(937);
CN_in_sigd(4005)	<=	VN_out_sigd(937);
CN_in_sigd(757)	<=	VN_out_sigd(938);
CN_in_sigd(2173)	<=	VN_out_sigd(938);
CN_in_sigd(3397)	<=	VN_out_sigd(938);
CN_in_sigd(4013)	<=	VN_out_sigd(938);
CN_in_sigd(765)	<=	VN_out_sigd(939);
CN_in_sigd(2181)	<=	VN_out_sigd(939);
CN_in_sigd(3405)	<=	VN_out_sigd(939);
CN_in_sigd(4021)	<=	VN_out_sigd(939);
CN_in_sigd(773)	<=	VN_out_sigd(940);
CN_in_sigd(2189)	<=	VN_out_sigd(940);
CN_in_sigd(3413)	<=	VN_out_sigd(940);
CN_in_sigd(4029)	<=	VN_out_sigd(940);
CN_in_sigd(781)	<=	VN_out_sigd(941);
CN_in_sigd(2197)	<=	VN_out_sigd(941);
CN_in_sigd(3421)	<=	VN_out_sigd(941);
CN_in_sigd(4037)	<=	VN_out_sigd(941);
CN_in_sigd(789)	<=	VN_out_sigd(942);
CN_in_sigd(2205)	<=	VN_out_sigd(942);
CN_in_sigd(3429)	<=	VN_out_sigd(942);
CN_in_sigd(4045)	<=	VN_out_sigd(942);
CN_in_sigd(797)	<=	VN_out_sigd(943);
CN_in_sigd(2213)	<=	VN_out_sigd(943);
CN_in_sigd(3437)	<=	VN_out_sigd(943);
CN_in_sigd(4053)	<=	VN_out_sigd(943);
CN_in_sigd(805)	<=	VN_out_sigd(944);
CN_in_sigd(2221)	<=	VN_out_sigd(944);
CN_in_sigd(3445)	<=	VN_out_sigd(944);
CN_in_sigd(4061)	<=	VN_out_sigd(944);
CN_in_sigd(813)	<=	VN_out_sigd(945);
CN_in_sigd(2229)	<=	VN_out_sigd(945);
CN_in_sigd(3453)	<=	VN_out_sigd(945);
CN_in_sigd(4069)	<=	VN_out_sigd(945);
CN_in_sigd(821)	<=	VN_out_sigd(946);
CN_in_sigd(2237)	<=	VN_out_sigd(946);
CN_in_sigd(3029)	<=	VN_out_sigd(946);
CN_in_sigd(4077)	<=	VN_out_sigd(946);
CN_in_sigd(829)	<=	VN_out_sigd(947);
CN_in_sigd(2245)	<=	VN_out_sigd(947);
CN_in_sigd(3037)	<=	VN_out_sigd(947);
CN_in_sigd(4085)	<=	VN_out_sigd(947);
CN_in_sigd(837)	<=	VN_out_sigd(948);
CN_in_sigd(2253)	<=	VN_out_sigd(948);
CN_in_sigd(3045)	<=	VN_out_sigd(948);
CN_in_sigd(4093)	<=	VN_out_sigd(948);
CN_in_sigd(845)	<=	VN_out_sigd(949);
CN_in_sigd(2261)	<=	VN_out_sigd(949);
CN_in_sigd(3053)	<=	VN_out_sigd(949);
CN_in_sigd(4101)	<=	VN_out_sigd(949);
CN_in_sigd(853)	<=	VN_out_sigd(950);
CN_in_sigd(2269)	<=	VN_out_sigd(950);
CN_in_sigd(3061)	<=	VN_out_sigd(950);
CN_in_sigd(4109)	<=	VN_out_sigd(950);
CN_in_sigd(861)	<=	VN_out_sigd(951);
CN_in_sigd(2277)	<=	VN_out_sigd(951);
CN_in_sigd(3069)	<=	VN_out_sigd(951);
CN_in_sigd(4117)	<=	VN_out_sigd(951);
CN_in_sigd(437)	<=	VN_out_sigd(952);
CN_in_sigd(2285)	<=	VN_out_sigd(952);
CN_in_sigd(3077)	<=	VN_out_sigd(952);
CN_in_sigd(4125)	<=	VN_out_sigd(952);
CN_in_sigd(445)	<=	VN_out_sigd(953);
CN_in_sigd(2293)	<=	VN_out_sigd(953);
CN_in_sigd(3085)	<=	VN_out_sigd(953);
CN_in_sigd(4133)	<=	VN_out_sigd(953);
CN_in_sigd(453)	<=	VN_out_sigd(954);
CN_in_sigd(2301)	<=	VN_out_sigd(954);
CN_in_sigd(3093)	<=	VN_out_sigd(954);
CN_in_sigd(4141)	<=	VN_out_sigd(954);
CN_in_sigd(461)	<=	VN_out_sigd(955);
CN_in_sigd(2309)	<=	VN_out_sigd(955);
CN_in_sigd(3101)	<=	VN_out_sigd(955);
CN_in_sigd(4149)	<=	VN_out_sigd(955);
CN_in_sigd(469)	<=	VN_out_sigd(956);
CN_in_sigd(2317)	<=	VN_out_sigd(956);
CN_in_sigd(3109)	<=	VN_out_sigd(956);
CN_in_sigd(4157)	<=	VN_out_sigd(956);
CN_in_sigd(477)	<=	VN_out_sigd(957);
CN_in_sigd(2325)	<=	VN_out_sigd(957);
CN_in_sigd(3117)	<=	VN_out_sigd(957);
CN_in_sigd(4165)	<=	VN_out_sigd(957);
CN_in_sigd(485)	<=	VN_out_sigd(958);
CN_in_sigd(2333)	<=	VN_out_sigd(958);
CN_in_sigd(3125)	<=	VN_out_sigd(958);
CN_in_sigd(4173)	<=	VN_out_sigd(958);
CN_in_sigd(493)	<=	VN_out_sigd(959);
CN_in_sigd(2341)	<=	VN_out_sigd(959);
CN_in_sigd(3133)	<=	VN_out_sigd(959);
CN_in_sigd(4181)	<=	VN_out_sigd(959);
CN_in_sigd(501)	<=	VN_out_sigd(960);
CN_in_sigd(2349)	<=	VN_out_sigd(960);
CN_in_sigd(3141)	<=	VN_out_sigd(960);
CN_in_sigd(4189)	<=	VN_out_sigd(960);
CN_in_sigd(509)	<=	VN_out_sigd(961);
CN_in_sigd(2357)	<=	VN_out_sigd(961);
CN_in_sigd(3149)	<=	VN_out_sigd(961);
CN_in_sigd(4197)	<=	VN_out_sigd(961);
CN_in_sigd(517)	<=	VN_out_sigd(962);
CN_in_sigd(2365)	<=	VN_out_sigd(962);
CN_in_sigd(3157)	<=	VN_out_sigd(962);
CN_in_sigd(4205)	<=	VN_out_sigd(962);
CN_in_sigd(525)	<=	VN_out_sigd(963);
CN_in_sigd(2373)	<=	VN_out_sigd(963);
CN_in_sigd(3165)	<=	VN_out_sigd(963);
CN_in_sigd(4213)	<=	VN_out_sigd(963);
CN_in_sigd(533)	<=	VN_out_sigd(964);
CN_in_sigd(2381)	<=	VN_out_sigd(964);
CN_in_sigd(3173)	<=	VN_out_sigd(964);
CN_in_sigd(4221)	<=	VN_out_sigd(964);
CN_in_sigd(541)	<=	VN_out_sigd(965);
CN_in_sigd(2389)	<=	VN_out_sigd(965);
CN_in_sigd(3181)	<=	VN_out_sigd(965);
CN_in_sigd(4229)	<=	VN_out_sigd(965);
CN_in_sigd(549)	<=	VN_out_sigd(966);
CN_in_sigd(2397)	<=	VN_out_sigd(966);
CN_in_sigd(3189)	<=	VN_out_sigd(966);
CN_in_sigd(4237)	<=	VN_out_sigd(966);
CN_in_sigd(557)	<=	VN_out_sigd(967);
CN_in_sigd(2405)	<=	VN_out_sigd(967);
CN_in_sigd(3197)	<=	VN_out_sigd(967);
CN_in_sigd(4245)	<=	VN_out_sigd(967);
CN_in_sigd(565)	<=	VN_out_sigd(968);
CN_in_sigd(2413)	<=	VN_out_sigd(968);
CN_in_sigd(3205)	<=	VN_out_sigd(968);
CN_in_sigd(4253)	<=	VN_out_sigd(968);
CN_in_sigd(573)	<=	VN_out_sigd(969);
CN_in_sigd(2421)	<=	VN_out_sigd(969);
CN_in_sigd(3213)	<=	VN_out_sigd(969);
CN_in_sigd(4261)	<=	VN_out_sigd(969);
CN_in_sigd(581)	<=	VN_out_sigd(970);
CN_in_sigd(2429)	<=	VN_out_sigd(970);
CN_in_sigd(3221)	<=	VN_out_sigd(970);
CN_in_sigd(4269)	<=	VN_out_sigd(970);
CN_in_sigd(589)	<=	VN_out_sigd(971);
CN_in_sigd(2437)	<=	VN_out_sigd(971);
CN_in_sigd(3229)	<=	VN_out_sigd(971);
CN_in_sigd(4277)	<=	VN_out_sigd(971);
CN_in_sigd(374)	<=	VN_out_sigd(972);
CN_in_sigd(1702)	<=	VN_out_sigd(972);
CN_in_sigd(3694)	<=	VN_out_sigd(972);
CN_in_sigd(5126)	<=	VN_out_sigd(972);
CN_in_sigd(382)	<=	VN_out_sigd(973);
CN_in_sigd(1710)	<=	VN_out_sigd(973);
CN_in_sigd(3702)	<=	VN_out_sigd(973);
CN_in_sigd(5134)	<=	VN_out_sigd(973);
CN_in_sigd(390)	<=	VN_out_sigd(974);
CN_in_sigd(1718)	<=	VN_out_sigd(974);
CN_in_sigd(3710)	<=	VN_out_sigd(974);
CN_in_sigd(5142)	<=	VN_out_sigd(974);
CN_in_sigd(398)	<=	VN_out_sigd(975);
CN_in_sigd(1726)	<=	VN_out_sigd(975);
CN_in_sigd(3718)	<=	VN_out_sigd(975);
CN_in_sigd(5150)	<=	VN_out_sigd(975);
CN_in_sigd(406)	<=	VN_out_sigd(976);
CN_in_sigd(1302)	<=	VN_out_sigd(976);
CN_in_sigd(3726)	<=	VN_out_sigd(976);
CN_in_sigd(5158)	<=	VN_out_sigd(976);
CN_in_sigd(414)	<=	VN_out_sigd(977);
CN_in_sigd(1310)	<=	VN_out_sigd(977);
CN_in_sigd(3734)	<=	VN_out_sigd(977);
CN_in_sigd(5166)	<=	VN_out_sigd(977);
CN_in_sigd(422)	<=	VN_out_sigd(978);
CN_in_sigd(1318)	<=	VN_out_sigd(978);
CN_in_sigd(3742)	<=	VN_out_sigd(978);
CN_in_sigd(5174)	<=	VN_out_sigd(978);
CN_in_sigd(430)	<=	VN_out_sigd(979);
CN_in_sigd(1326)	<=	VN_out_sigd(979);
CN_in_sigd(3750)	<=	VN_out_sigd(979);
CN_in_sigd(5182)	<=	VN_out_sigd(979);
CN_in_sigd(6)	<=	VN_out_sigd(980);
CN_in_sigd(1334)	<=	VN_out_sigd(980);
CN_in_sigd(3758)	<=	VN_out_sigd(980);
CN_in_sigd(4758)	<=	VN_out_sigd(980);
CN_in_sigd(14)	<=	VN_out_sigd(981);
CN_in_sigd(1342)	<=	VN_out_sigd(981);
CN_in_sigd(3766)	<=	VN_out_sigd(981);
CN_in_sigd(4766)	<=	VN_out_sigd(981);
CN_in_sigd(22)	<=	VN_out_sigd(982);
CN_in_sigd(1350)	<=	VN_out_sigd(982);
CN_in_sigd(3774)	<=	VN_out_sigd(982);
CN_in_sigd(4774)	<=	VN_out_sigd(982);
CN_in_sigd(30)	<=	VN_out_sigd(983);
CN_in_sigd(1358)	<=	VN_out_sigd(983);
CN_in_sigd(3782)	<=	VN_out_sigd(983);
CN_in_sigd(4782)	<=	VN_out_sigd(983);
CN_in_sigd(38)	<=	VN_out_sigd(984);
CN_in_sigd(1366)	<=	VN_out_sigd(984);
CN_in_sigd(3790)	<=	VN_out_sigd(984);
CN_in_sigd(4790)	<=	VN_out_sigd(984);
CN_in_sigd(46)	<=	VN_out_sigd(985);
CN_in_sigd(1374)	<=	VN_out_sigd(985);
CN_in_sigd(3798)	<=	VN_out_sigd(985);
CN_in_sigd(4798)	<=	VN_out_sigd(985);
CN_in_sigd(54)	<=	VN_out_sigd(986);
CN_in_sigd(1382)	<=	VN_out_sigd(986);
CN_in_sigd(3806)	<=	VN_out_sigd(986);
CN_in_sigd(4806)	<=	VN_out_sigd(986);
CN_in_sigd(62)	<=	VN_out_sigd(987);
CN_in_sigd(1390)	<=	VN_out_sigd(987);
CN_in_sigd(3814)	<=	VN_out_sigd(987);
CN_in_sigd(4814)	<=	VN_out_sigd(987);
CN_in_sigd(70)	<=	VN_out_sigd(988);
CN_in_sigd(1398)	<=	VN_out_sigd(988);
CN_in_sigd(3822)	<=	VN_out_sigd(988);
CN_in_sigd(4822)	<=	VN_out_sigd(988);
CN_in_sigd(78)	<=	VN_out_sigd(989);
CN_in_sigd(1406)	<=	VN_out_sigd(989);
CN_in_sigd(3830)	<=	VN_out_sigd(989);
CN_in_sigd(4830)	<=	VN_out_sigd(989);
CN_in_sigd(86)	<=	VN_out_sigd(990);
CN_in_sigd(1414)	<=	VN_out_sigd(990);
CN_in_sigd(3838)	<=	VN_out_sigd(990);
CN_in_sigd(4838)	<=	VN_out_sigd(990);
CN_in_sigd(94)	<=	VN_out_sigd(991);
CN_in_sigd(1422)	<=	VN_out_sigd(991);
CN_in_sigd(3846)	<=	VN_out_sigd(991);
CN_in_sigd(4846)	<=	VN_out_sigd(991);
CN_in_sigd(102)	<=	VN_out_sigd(992);
CN_in_sigd(1430)	<=	VN_out_sigd(992);
CN_in_sigd(3854)	<=	VN_out_sigd(992);
CN_in_sigd(4854)	<=	VN_out_sigd(992);
CN_in_sigd(110)	<=	VN_out_sigd(993);
CN_in_sigd(1438)	<=	VN_out_sigd(993);
CN_in_sigd(3862)	<=	VN_out_sigd(993);
CN_in_sigd(4862)	<=	VN_out_sigd(993);
CN_in_sigd(118)	<=	VN_out_sigd(994);
CN_in_sigd(1446)	<=	VN_out_sigd(994);
CN_in_sigd(3870)	<=	VN_out_sigd(994);
CN_in_sigd(4870)	<=	VN_out_sigd(994);
CN_in_sigd(126)	<=	VN_out_sigd(995);
CN_in_sigd(1454)	<=	VN_out_sigd(995);
CN_in_sigd(3878)	<=	VN_out_sigd(995);
CN_in_sigd(4878)	<=	VN_out_sigd(995);
CN_in_sigd(134)	<=	VN_out_sigd(996);
CN_in_sigd(1462)	<=	VN_out_sigd(996);
CN_in_sigd(3886)	<=	VN_out_sigd(996);
CN_in_sigd(4886)	<=	VN_out_sigd(996);
CN_in_sigd(142)	<=	VN_out_sigd(997);
CN_in_sigd(1470)	<=	VN_out_sigd(997);
CN_in_sigd(3462)	<=	VN_out_sigd(997);
CN_in_sigd(4894)	<=	VN_out_sigd(997);
CN_in_sigd(150)	<=	VN_out_sigd(998);
CN_in_sigd(1478)	<=	VN_out_sigd(998);
CN_in_sigd(3470)	<=	VN_out_sigd(998);
CN_in_sigd(4902)	<=	VN_out_sigd(998);
CN_in_sigd(158)	<=	VN_out_sigd(999);
CN_in_sigd(1486)	<=	VN_out_sigd(999);
CN_in_sigd(3478)	<=	VN_out_sigd(999);
CN_in_sigd(4910)	<=	VN_out_sigd(999);
CN_in_sigd(166)	<=	VN_out_sigd(1000);
CN_in_sigd(1494)	<=	VN_out_sigd(1000);
CN_in_sigd(3486)	<=	VN_out_sigd(1000);
CN_in_sigd(4918)	<=	VN_out_sigd(1000);
CN_in_sigd(174)	<=	VN_out_sigd(1001);
CN_in_sigd(1502)	<=	VN_out_sigd(1001);
CN_in_sigd(3494)	<=	VN_out_sigd(1001);
CN_in_sigd(4926)	<=	VN_out_sigd(1001);
CN_in_sigd(182)	<=	VN_out_sigd(1002);
CN_in_sigd(1510)	<=	VN_out_sigd(1002);
CN_in_sigd(3502)	<=	VN_out_sigd(1002);
CN_in_sigd(4934)	<=	VN_out_sigd(1002);
CN_in_sigd(190)	<=	VN_out_sigd(1003);
CN_in_sigd(1518)	<=	VN_out_sigd(1003);
CN_in_sigd(3510)	<=	VN_out_sigd(1003);
CN_in_sigd(4942)	<=	VN_out_sigd(1003);
CN_in_sigd(198)	<=	VN_out_sigd(1004);
CN_in_sigd(1526)	<=	VN_out_sigd(1004);
CN_in_sigd(3518)	<=	VN_out_sigd(1004);
CN_in_sigd(4950)	<=	VN_out_sigd(1004);
CN_in_sigd(206)	<=	VN_out_sigd(1005);
CN_in_sigd(1534)	<=	VN_out_sigd(1005);
CN_in_sigd(3526)	<=	VN_out_sigd(1005);
CN_in_sigd(4958)	<=	VN_out_sigd(1005);
CN_in_sigd(214)	<=	VN_out_sigd(1006);
CN_in_sigd(1542)	<=	VN_out_sigd(1006);
CN_in_sigd(3534)	<=	VN_out_sigd(1006);
CN_in_sigd(4966)	<=	VN_out_sigd(1006);
CN_in_sigd(222)	<=	VN_out_sigd(1007);
CN_in_sigd(1550)	<=	VN_out_sigd(1007);
CN_in_sigd(3542)	<=	VN_out_sigd(1007);
CN_in_sigd(4974)	<=	VN_out_sigd(1007);
CN_in_sigd(230)	<=	VN_out_sigd(1008);
CN_in_sigd(1558)	<=	VN_out_sigd(1008);
CN_in_sigd(3550)	<=	VN_out_sigd(1008);
CN_in_sigd(4982)	<=	VN_out_sigd(1008);
CN_in_sigd(238)	<=	VN_out_sigd(1009);
CN_in_sigd(1566)	<=	VN_out_sigd(1009);
CN_in_sigd(3558)	<=	VN_out_sigd(1009);
CN_in_sigd(4990)	<=	VN_out_sigd(1009);
CN_in_sigd(246)	<=	VN_out_sigd(1010);
CN_in_sigd(1574)	<=	VN_out_sigd(1010);
CN_in_sigd(3566)	<=	VN_out_sigd(1010);
CN_in_sigd(4998)	<=	VN_out_sigd(1010);
CN_in_sigd(254)	<=	VN_out_sigd(1011);
CN_in_sigd(1582)	<=	VN_out_sigd(1011);
CN_in_sigd(3574)	<=	VN_out_sigd(1011);
CN_in_sigd(5006)	<=	VN_out_sigd(1011);
CN_in_sigd(262)	<=	VN_out_sigd(1012);
CN_in_sigd(1590)	<=	VN_out_sigd(1012);
CN_in_sigd(3582)	<=	VN_out_sigd(1012);
CN_in_sigd(5014)	<=	VN_out_sigd(1012);
CN_in_sigd(270)	<=	VN_out_sigd(1013);
CN_in_sigd(1598)	<=	VN_out_sigd(1013);
CN_in_sigd(3590)	<=	VN_out_sigd(1013);
CN_in_sigd(5022)	<=	VN_out_sigd(1013);
CN_in_sigd(278)	<=	VN_out_sigd(1014);
CN_in_sigd(1606)	<=	VN_out_sigd(1014);
CN_in_sigd(3598)	<=	VN_out_sigd(1014);
CN_in_sigd(5030)	<=	VN_out_sigd(1014);
CN_in_sigd(286)	<=	VN_out_sigd(1015);
CN_in_sigd(1614)	<=	VN_out_sigd(1015);
CN_in_sigd(3606)	<=	VN_out_sigd(1015);
CN_in_sigd(5038)	<=	VN_out_sigd(1015);
CN_in_sigd(294)	<=	VN_out_sigd(1016);
CN_in_sigd(1622)	<=	VN_out_sigd(1016);
CN_in_sigd(3614)	<=	VN_out_sigd(1016);
CN_in_sigd(5046)	<=	VN_out_sigd(1016);
CN_in_sigd(302)	<=	VN_out_sigd(1017);
CN_in_sigd(1630)	<=	VN_out_sigd(1017);
CN_in_sigd(3622)	<=	VN_out_sigd(1017);
CN_in_sigd(5054)	<=	VN_out_sigd(1017);
CN_in_sigd(310)	<=	VN_out_sigd(1018);
CN_in_sigd(1638)	<=	VN_out_sigd(1018);
CN_in_sigd(3630)	<=	VN_out_sigd(1018);
CN_in_sigd(5062)	<=	VN_out_sigd(1018);
CN_in_sigd(318)	<=	VN_out_sigd(1019);
CN_in_sigd(1646)	<=	VN_out_sigd(1019);
CN_in_sigd(3638)	<=	VN_out_sigd(1019);
CN_in_sigd(5070)	<=	VN_out_sigd(1019);
CN_in_sigd(326)	<=	VN_out_sigd(1020);
CN_in_sigd(1654)	<=	VN_out_sigd(1020);
CN_in_sigd(3646)	<=	VN_out_sigd(1020);
CN_in_sigd(5078)	<=	VN_out_sigd(1020);
CN_in_sigd(334)	<=	VN_out_sigd(1021);
CN_in_sigd(1662)	<=	VN_out_sigd(1021);
CN_in_sigd(3654)	<=	VN_out_sigd(1021);
CN_in_sigd(5086)	<=	VN_out_sigd(1021);
CN_in_sigd(342)	<=	VN_out_sigd(1022);
CN_in_sigd(1670)	<=	VN_out_sigd(1022);
CN_in_sigd(3662)	<=	VN_out_sigd(1022);
CN_in_sigd(5094)	<=	VN_out_sigd(1022);
CN_in_sigd(350)	<=	VN_out_sigd(1023);
CN_in_sigd(1678)	<=	VN_out_sigd(1023);
CN_in_sigd(3670)	<=	VN_out_sigd(1023);
CN_in_sigd(5102)	<=	VN_out_sigd(1023);
CN_in_sigd(358)	<=	VN_out_sigd(1024);
CN_in_sigd(1686)	<=	VN_out_sigd(1024);
CN_in_sigd(3678)	<=	VN_out_sigd(1024);
CN_in_sigd(5110)	<=	VN_out_sigd(1024);
CN_in_sigd(366)	<=	VN_out_sigd(1025);
CN_in_sigd(1694)	<=	VN_out_sigd(1025);
CN_in_sigd(3686)	<=	VN_out_sigd(1025);
CN_in_sigd(5118)	<=	VN_out_sigd(1025);
CN_in_sigd(750)	<=	VN_out_sigd(1026);
CN_in_sigd(2294)	<=	VN_out_sigd(1026);
CN_in_sigd(2694)	<=	VN_out_sigd(1026);
CN_in_sigd(4046)	<=	VN_out_sigd(1026);
CN_in_sigd(758)	<=	VN_out_sigd(1027);
CN_in_sigd(2302)	<=	VN_out_sigd(1027);
CN_in_sigd(2702)	<=	VN_out_sigd(1027);
CN_in_sigd(4054)	<=	VN_out_sigd(1027);
CN_in_sigd(766)	<=	VN_out_sigd(1028);
CN_in_sigd(2310)	<=	VN_out_sigd(1028);
CN_in_sigd(2710)	<=	VN_out_sigd(1028);
CN_in_sigd(4062)	<=	VN_out_sigd(1028);
CN_in_sigd(774)	<=	VN_out_sigd(1029);
CN_in_sigd(2318)	<=	VN_out_sigd(1029);
CN_in_sigd(2718)	<=	VN_out_sigd(1029);
CN_in_sigd(4070)	<=	VN_out_sigd(1029);
CN_in_sigd(782)	<=	VN_out_sigd(1030);
CN_in_sigd(2326)	<=	VN_out_sigd(1030);
CN_in_sigd(2726)	<=	VN_out_sigd(1030);
CN_in_sigd(4078)	<=	VN_out_sigd(1030);
CN_in_sigd(790)	<=	VN_out_sigd(1031);
CN_in_sigd(2334)	<=	VN_out_sigd(1031);
CN_in_sigd(2734)	<=	VN_out_sigd(1031);
CN_in_sigd(4086)	<=	VN_out_sigd(1031);
CN_in_sigd(798)	<=	VN_out_sigd(1032);
CN_in_sigd(2342)	<=	VN_out_sigd(1032);
CN_in_sigd(2742)	<=	VN_out_sigd(1032);
CN_in_sigd(4094)	<=	VN_out_sigd(1032);
CN_in_sigd(806)	<=	VN_out_sigd(1033);
CN_in_sigd(2350)	<=	VN_out_sigd(1033);
CN_in_sigd(2750)	<=	VN_out_sigd(1033);
CN_in_sigd(4102)	<=	VN_out_sigd(1033);
CN_in_sigd(814)	<=	VN_out_sigd(1034);
CN_in_sigd(2358)	<=	VN_out_sigd(1034);
CN_in_sigd(2758)	<=	VN_out_sigd(1034);
CN_in_sigd(4110)	<=	VN_out_sigd(1034);
CN_in_sigd(822)	<=	VN_out_sigd(1035);
CN_in_sigd(2366)	<=	VN_out_sigd(1035);
CN_in_sigd(2766)	<=	VN_out_sigd(1035);
CN_in_sigd(4118)	<=	VN_out_sigd(1035);
CN_in_sigd(830)	<=	VN_out_sigd(1036);
CN_in_sigd(2374)	<=	VN_out_sigd(1036);
CN_in_sigd(2774)	<=	VN_out_sigd(1036);
CN_in_sigd(4126)	<=	VN_out_sigd(1036);
CN_in_sigd(838)	<=	VN_out_sigd(1037);
CN_in_sigd(2382)	<=	VN_out_sigd(1037);
CN_in_sigd(2782)	<=	VN_out_sigd(1037);
CN_in_sigd(4134)	<=	VN_out_sigd(1037);
CN_in_sigd(846)	<=	VN_out_sigd(1038);
CN_in_sigd(2390)	<=	VN_out_sigd(1038);
CN_in_sigd(2790)	<=	VN_out_sigd(1038);
CN_in_sigd(4142)	<=	VN_out_sigd(1038);
CN_in_sigd(854)	<=	VN_out_sigd(1039);
CN_in_sigd(2398)	<=	VN_out_sigd(1039);
CN_in_sigd(2798)	<=	VN_out_sigd(1039);
CN_in_sigd(4150)	<=	VN_out_sigd(1039);
CN_in_sigd(862)	<=	VN_out_sigd(1040);
CN_in_sigd(2406)	<=	VN_out_sigd(1040);
CN_in_sigd(2806)	<=	VN_out_sigd(1040);
CN_in_sigd(4158)	<=	VN_out_sigd(1040);
CN_in_sigd(438)	<=	VN_out_sigd(1041);
CN_in_sigd(2414)	<=	VN_out_sigd(1041);
CN_in_sigd(2814)	<=	VN_out_sigd(1041);
CN_in_sigd(4166)	<=	VN_out_sigd(1041);
CN_in_sigd(446)	<=	VN_out_sigd(1042);
CN_in_sigd(2422)	<=	VN_out_sigd(1042);
CN_in_sigd(2822)	<=	VN_out_sigd(1042);
CN_in_sigd(4174)	<=	VN_out_sigd(1042);
CN_in_sigd(454)	<=	VN_out_sigd(1043);
CN_in_sigd(2430)	<=	VN_out_sigd(1043);
CN_in_sigd(2830)	<=	VN_out_sigd(1043);
CN_in_sigd(4182)	<=	VN_out_sigd(1043);
CN_in_sigd(462)	<=	VN_out_sigd(1044);
CN_in_sigd(2438)	<=	VN_out_sigd(1044);
CN_in_sigd(2838)	<=	VN_out_sigd(1044);
CN_in_sigd(4190)	<=	VN_out_sigd(1044);
CN_in_sigd(470)	<=	VN_out_sigd(1045);
CN_in_sigd(2446)	<=	VN_out_sigd(1045);
CN_in_sigd(2846)	<=	VN_out_sigd(1045);
CN_in_sigd(4198)	<=	VN_out_sigd(1045);
CN_in_sigd(478)	<=	VN_out_sigd(1046);
CN_in_sigd(2454)	<=	VN_out_sigd(1046);
CN_in_sigd(2854)	<=	VN_out_sigd(1046);
CN_in_sigd(4206)	<=	VN_out_sigd(1046);
CN_in_sigd(486)	<=	VN_out_sigd(1047);
CN_in_sigd(2462)	<=	VN_out_sigd(1047);
CN_in_sigd(2862)	<=	VN_out_sigd(1047);
CN_in_sigd(4214)	<=	VN_out_sigd(1047);
CN_in_sigd(494)	<=	VN_out_sigd(1048);
CN_in_sigd(2470)	<=	VN_out_sigd(1048);
CN_in_sigd(2870)	<=	VN_out_sigd(1048);
CN_in_sigd(4222)	<=	VN_out_sigd(1048);
CN_in_sigd(502)	<=	VN_out_sigd(1049);
CN_in_sigd(2478)	<=	VN_out_sigd(1049);
CN_in_sigd(2878)	<=	VN_out_sigd(1049);
CN_in_sigd(4230)	<=	VN_out_sigd(1049);
CN_in_sigd(510)	<=	VN_out_sigd(1050);
CN_in_sigd(2486)	<=	VN_out_sigd(1050);
CN_in_sigd(2886)	<=	VN_out_sigd(1050);
CN_in_sigd(4238)	<=	VN_out_sigd(1050);
CN_in_sigd(518)	<=	VN_out_sigd(1051);
CN_in_sigd(2494)	<=	VN_out_sigd(1051);
CN_in_sigd(2894)	<=	VN_out_sigd(1051);
CN_in_sigd(4246)	<=	VN_out_sigd(1051);
CN_in_sigd(526)	<=	VN_out_sigd(1052);
CN_in_sigd(2502)	<=	VN_out_sigd(1052);
CN_in_sigd(2902)	<=	VN_out_sigd(1052);
CN_in_sigd(4254)	<=	VN_out_sigd(1052);
CN_in_sigd(534)	<=	VN_out_sigd(1053);
CN_in_sigd(2510)	<=	VN_out_sigd(1053);
CN_in_sigd(2910)	<=	VN_out_sigd(1053);
CN_in_sigd(4262)	<=	VN_out_sigd(1053);
CN_in_sigd(542)	<=	VN_out_sigd(1054);
CN_in_sigd(2518)	<=	VN_out_sigd(1054);
CN_in_sigd(2918)	<=	VN_out_sigd(1054);
CN_in_sigd(4270)	<=	VN_out_sigd(1054);
CN_in_sigd(550)	<=	VN_out_sigd(1055);
CN_in_sigd(2526)	<=	VN_out_sigd(1055);
CN_in_sigd(2926)	<=	VN_out_sigd(1055);
CN_in_sigd(4278)	<=	VN_out_sigd(1055);
CN_in_sigd(558)	<=	VN_out_sigd(1056);
CN_in_sigd(2534)	<=	VN_out_sigd(1056);
CN_in_sigd(2934)	<=	VN_out_sigd(1056);
CN_in_sigd(4286)	<=	VN_out_sigd(1056);
CN_in_sigd(566)	<=	VN_out_sigd(1057);
CN_in_sigd(2542)	<=	VN_out_sigd(1057);
CN_in_sigd(2942)	<=	VN_out_sigd(1057);
CN_in_sigd(4294)	<=	VN_out_sigd(1057);
CN_in_sigd(574)	<=	VN_out_sigd(1058);
CN_in_sigd(2550)	<=	VN_out_sigd(1058);
CN_in_sigd(2950)	<=	VN_out_sigd(1058);
CN_in_sigd(4302)	<=	VN_out_sigd(1058);
CN_in_sigd(582)	<=	VN_out_sigd(1059);
CN_in_sigd(2558)	<=	VN_out_sigd(1059);
CN_in_sigd(2958)	<=	VN_out_sigd(1059);
CN_in_sigd(4310)	<=	VN_out_sigd(1059);
CN_in_sigd(590)	<=	VN_out_sigd(1060);
CN_in_sigd(2566)	<=	VN_out_sigd(1060);
CN_in_sigd(2966)	<=	VN_out_sigd(1060);
CN_in_sigd(4318)	<=	VN_out_sigd(1060);
CN_in_sigd(598)	<=	VN_out_sigd(1061);
CN_in_sigd(2574)	<=	VN_out_sigd(1061);
CN_in_sigd(2974)	<=	VN_out_sigd(1061);
CN_in_sigd(3894)	<=	VN_out_sigd(1061);
CN_in_sigd(606)	<=	VN_out_sigd(1062);
CN_in_sigd(2582)	<=	VN_out_sigd(1062);
CN_in_sigd(2982)	<=	VN_out_sigd(1062);
CN_in_sigd(3902)	<=	VN_out_sigd(1062);
CN_in_sigd(614)	<=	VN_out_sigd(1063);
CN_in_sigd(2590)	<=	VN_out_sigd(1063);
CN_in_sigd(2990)	<=	VN_out_sigd(1063);
CN_in_sigd(3910)	<=	VN_out_sigd(1063);
CN_in_sigd(622)	<=	VN_out_sigd(1064);
CN_in_sigd(2166)	<=	VN_out_sigd(1064);
CN_in_sigd(2998)	<=	VN_out_sigd(1064);
CN_in_sigd(3918)	<=	VN_out_sigd(1064);
CN_in_sigd(630)	<=	VN_out_sigd(1065);
CN_in_sigd(2174)	<=	VN_out_sigd(1065);
CN_in_sigd(3006)	<=	VN_out_sigd(1065);
CN_in_sigd(3926)	<=	VN_out_sigd(1065);
CN_in_sigd(638)	<=	VN_out_sigd(1066);
CN_in_sigd(2182)	<=	VN_out_sigd(1066);
CN_in_sigd(3014)	<=	VN_out_sigd(1066);
CN_in_sigd(3934)	<=	VN_out_sigd(1066);
CN_in_sigd(646)	<=	VN_out_sigd(1067);
CN_in_sigd(2190)	<=	VN_out_sigd(1067);
CN_in_sigd(3022)	<=	VN_out_sigd(1067);
CN_in_sigd(3942)	<=	VN_out_sigd(1067);
CN_in_sigd(654)	<=	VN_out_sigd(1068);
CN_in_sigd(2198)	<=	VN_out_sigd(1068);
CN_in_sigd(2598)	<=	VN_out_sigd(1068);
CN_in_sigd(3950)	<=	VN_out_sigd(1068);
CN_in_sigd(662)	<=	VN_out_sigd(1069);
CN_in_sigd(2206)	<=	VN_out_sigd(1069);
CN_in_sigd(2606)	<=	VN_out_sigd(1069);
CN_in_sigd(3958)	<=	VN_out_sigd(1069);
CN_in_sigd(670)	<=	VN_out_sigd(1070);
CN_in_sigd(2214)	<=	VN_out_sigd(1070);
CN_in_sigd(2614)	<=	VN_out_sigd(1070);
CN_in_sigd(3966)	<=	VN_out_sigd(1070);
CN_in_sigd(678)	<=	VN_out_sigd(1071);
CN_in_sigd(2222)	<=	VN_out_sigd(1071);
CN_in_sigd(2622)	<=	VN_out_sigd(1071);
CN_in_sigd(3974)	<=	VN_out_sigd(1071);
CN_in_sigd(686)	<=	VN_out_sigd(1072);
CN_in_sigd(2230)	<=	VN_out_sigd(1072);
CN_in_sigd(2630)	<=	VN_out_sigd(1072);
CN_in_sigd(3982)	<=	VN_out_sigd(1072);
CN_in_sigd(694)	<=	VN_out_sigd(1073);
CN_in_sigd(2238)	<=	VN_out_sigd(1073);
CN_in_sigd(2638)	<=	VN_out_sigd(1073);
CN_in_sigd(3990)	<=	VN_out_sigd(1073);
CN_in_sigd(702)	<=	VN_out_sigd(1074);
CN_in_sigd(2246)	<=	VN_out_sigd(1074);
CN_in_sigd(2646)	<=	VN_out_sigd(1074);
CN_in_sigd(3998)	<=	VN_out_sigd(1074);
CN_in_sigd(710)	<=	VN_out_sigd(1075);
CN_in_sigd(2254)	<=	VN_out_sigd(1075);
CN_in_sigd(2654)	<=	VN_out_sigd(1075);
CN_in_sigd(4006)	<=	VN_out_sigd(1075);
CN_in_sigd(718)	<=	VN_out_sigd(1076);
CN_in_sigd(2262)	<=	VN_out_sigd(1076);
CN_in_sigd(2662)	<=	VN_out_sigd(1076);
CN_in_sigd(4014)	<=	VN_out_sigd(1076);
CN_in_sigd(726)	<=	VN_out_sigd(1077);
CN_in_sigd(2270)	<=	VN_out_sigd(1077);
CN_in_sigd(2670)	<=	VN_out_sigd(1077);
CN_in_sigd(4022)	<=	VN_out_sigd(1077);
CN_in_sigd(734)	<=	VN_out_sigd(1078);
CN_in_sigd(2278)	<=	VN_out_sigd(1078);
CN_in_sigd(2678)	<=	VN_out_sigd(1078);
CN_in_sigd(4030)	<=	VN_out_sigd(1078);
CN_in_sigd(742)	<=	VN_out_sigd(1079);
CN_in_sigd(2286)	<=	VN_out_sigd(1079);
CN_in_sigd(2686)	<=	VN_out_sigd(1079);
CN_in_sigd(4038)	<=	VN_out_sigd(1079);
CN_in_sigd(1062)	<=	VN_out_sigd(1080);
CN_in_sigd(1806)	<=	VN_out_sigd(1080);
CN_in_sigd(3238)	<=	VN_out_sigd(1080);
CN_in_sigd(4470)	<=	VN_out_sigd(1080);
CN_in_sigd(1070)	<=	VN_out_sigd(1081);
CN_in_sigd(1814)	<=	VN_out_sigd(1081);
CN_in_sigd(3246)	<=	VN_out_sigd(1081);
CN_in_sigd(4478)	<=	VN_out_sigd(1081);
CN_in_sigd(1078)	<=	VN_out_sigd(1082);
CN_in_sigd(1822)	<=	VN_out_sigd(1082);
CN_in_sigd(3254)	<=	VN_out_sigd(1082);
CN_in_sigd(4486)	<=	VN_out_sigd(1082);
CN_in_sigd(1086)	<=	VN_out_sigd(1083);
CN_in_sigd(1830)	<=	VN_out_sigd(1083);
CN_in_sigd(3262)	<=	VN_out_sigd(1083);
CN_in_sigd(4494)	<=	VN_out_sigd(1083);
CN_in_sigd(1094)	<=	VN_out_sigd(1084);
CN_in_sigd(1838)	<=	VN_out_sigd(1084);
CN_in_sigd(3270)	<=	VN_out_sigd(1084);
CN_in_sigd(4502)	<=	VN_out_sigd(1084);
CN_in_sigd(1102)	<=	VN_out_sigd(1085);
CN_in_sigd(1846)	<=	VN_out_sigd(1085);
CN_in_sigd(3278)	<=	VN_out_sigd(1085);
CN_in_sigd(4510)	<=	VN_out_sigd(1085);
CN_in_sigd(1110)	<=	VN_out_sigd(1086);
CN_in_sigd(1854)	<=	VN_out_sigd(1086);
CN_in_sigd(3286)	<=	VN_out_sigd(1086);
CN_in_sigd(4518)	<=	VN_out_sigd(1086);
CN_in_sigd(1118)	<=	VN_out_sigd(1087);
CN_in_sigd(1862)	<=	VN_out_sigd(1087);
CN_in_sigd(3294)	<=	VN_out_sigd(1087);
CN_in_sigd(4526)	<=	VN_out_sigd(1087);
CN_in_sigd(1126)	<=	VN_out_sigd(1088);
CN_in_sigd(1870)	<=	VN_out_sigd(1088);
CN_in_sigd(3302)	<=	VN_out_sigd(1088);
CN_in_sigd(4534)	<=	VN_out_sigd(1088);
CN_in_sigd(1134)	<=	VN_out_sigd(1089);
CN_in_sigd(1878)	<=	VN_out_sigd(1089);
CN_in_sigd(3310)	<=	VN_out_sigd(1089);
CN_in_sigd(4542)	<=	VN_out_sigd(1089);
CN_in_sigd(1142)	<=	VN_out_sigd(1090);
CN_in_sigd(1886)	<=	VN_out_sigd(1090);
CN_in_sigd(3318)	<=	VN_out_sigd(1090);
CN_in_sigd(4550)	<=	VN_out_sigd(1090);
CN_in_sigd(1150)	<=	VN_out_sigd(1091);
CN_in_sigd(1894)	<=	VN_out_sigd(1091);
CN_in_sigd(3326)	<=	VN_out_sigd(1091);
CN_in_sigd(4558)	<=	VN_out_sigd(1091);
CN_in_sigd(1158)	<=	VN_out_sigd(1092);
CN_in_sigd(1902)	<=	VN_out_sigd(1092);
CN_in_sigd(3334)	<=	VN_out_sigd(1092);
CN_in_sigd(4566)	<=	VN_out_sigd(1092);
CN_in_sigd(1166)	<=	VN_out_sigd(1093);
CN_in_sigd(1910)	<=	VN_out_sigd(1093);
CN_in_sigd(3342)	<=	VN_out_sigd(1093);
CN_in_sigd(4574)	<=	VN_out_sigd(1093);
CN_in_sigd(1174)	<=	VN_out_sigd(1094);
CN_in_sigd(1918)	<=	VN_out_sigd(1094);
CN_in_sigd(3350)	<=	VN_out_sigd(1094);
CN_in_sigd(4582)	<=	VN_out_sigd(1094);
CN_in_sigd(1182)	<=	VN_out_sigd(1095);
CN_in_sigd(1926)	<=	VN_out_sigd(1095);
CN_in_sigd(3358)	<=	VN_out_sigd(1095);
CN_in_sigd(4590)	<=	VN_out_sigd(1095);
CN_in_sigd(1190)	<=	VN_out_sigd(1096);
CN_in_sigd(1934)	<=	VN_out_sigd(1096);
CN_in_sigd(3366)	<=	VN_out_sigd(1096);
CN_in_sigd(4598)	<=	VN_out_sigd(1096);
CN_in_sigd(1198)	<=	VN_out_sigd(1097);
CN_in_sigd(1942)	<=	VN_out_sigd(1097);
CN_in_sigd(3374)	<=	VN_out_sigd(1097);
CN_in_sigd(4606)	<=	VN_out_sigd(1097);
CN_in_sigd(1206)	<=	VN_out_sigd(1098);
CN_in_sigd(1950)	<=	VN_out_sigd(1098);
CN_in_sigd(3382)	<=	VN_out_sigd(1098);
CN_in_sigd(4614)	<=	VN_out_sigd(1098);
CN_in_sigd(1214)	<=	VN_out_sigd(1099);
CN_in_sigd(1958)	<=	VN_out_sigd(1099);
CN_in_sigd(3390)	<=	VN_out_sigd(1099);
CN_in_sigd(4622)	<=	VN_out_sigd(1099);
CN_in_sigd(1222)	<=	VN_out_sigd(1100);
CN_in_sigd(1966)	<=	VN_out_sigd(1100);
CN_in_sigd(3398)	<=	VN_out_sigd(1100);
CN_in_sigd(4630)	<=	VN_out_sigd(1100);
CN_in_sigd(1230)	<=	VN_out_sigd(1101);
CN_in_sigd(1974)	<=	VN_out_sigd(1101);
CN_in_sigd(3406)	<=	VN_out_sigd(1101);
CN_in_sigd(4638)	<=	VN_out_sigd(1101);
CN_in_sigd(1238)	<=	VN_out_sigd(1102);
CN_in_sigd(1982)	<=	VN_out_sigd(1102);
CN_in_sigd(3414)	<=	VN_out_sigd(1102);
CN_in_sigd(4646)	<=	VN_out_sigd(1102);
CN_in_sigd(1246)	<=	VN_out_sigd(1103);
CN_in_sigd(1990)	<=	VN_out_sigd(1103);
CN_in_sigd(3422)	<=	VN_out_sigd(1103);
CN_in_sigd(4654)	<=	VN_out_sigd(1103);
CN_in_sigd(1254)	<=	VN_out_sigd(1104);
CN_in_sigd(1998)	<=	VN_out_sigd(1104);
CN_in_sigd(3430)	<=	VN_out_sigd(1104);
CN_in_sigd(4662)	<=	VN_out_sigd(1104);
CN_in_sigd(1262)	<=	VN_out_sigd(1105);
CN_in_sigd(2006)	<=	VN_out_sigd(1105);
CN_in_sigd(3438)	<=	VN_out_sigd(1105);
CN_in_sigd(4670)	<=	VN_out_sigd(1105);
CN_in_sigd(1270)	<=	VN_out_sigd(1106);
CN_in_sigd(2014)	<=	VN_out_sigd(1106);
CN_in_sigd(3446)	<=	VN_out_sigd(1106);
CN_in_sigd(4678)	<=	VN_out_sigd(1106);
CN_in_sigd(1278)	<=	VN_out_sigd(1107);
CN_in_sigd(2022)	<=	VN_out_sigd(1107);
CN_in_sigd(3454)	<=	VN_out_sigd(1107);
CN_in_sigd(4686)	<=	VN_out_sigd(1107);
CN_in_sigd(1286)	<=	VN_out_sigd(1108);
CN_in_sigd(2030)	<=	VN_out_sigd(1108);
CN_in_sigd(3030)	<=	VN_out_sigd(1108);
CN_in_sigd(4694)	<=	VN_out_sigd(1108);
CN_in_sigd(1294)	<=	VN_out_sigd(1109);
CN_in_sigd(2038)	<=	VN_out_sigd(1109);
CN_in_sigd(3038)	<=	VN_out_sigd(1109);
CN_in_sigd(4702)	<=	VN_out_sigd(1109);
CN_in_sigd(870)	<=	VN_out_sigd(1110);
CN_in_sigd(2046)	<=	VN_out_sigd(1110);
CN_in_sigd(3046)	<=	VN_out_sigd(1110);
CN_in_sigd(4710)	<=	VN_out_sigd(1110);
CN_in_sigd(878)	<=	VN_out_sigd(1111);
CN_in_sigd(2054)	<=	VN_out_sigd(1111);
CN_in_sigd(3054)	<=	VN_out_sigd(1111);
CN_in_sigd(4718)	<=	VN_out_sigd(1111);
CN_in_sigd(886)	<=	VN_out_sigd(1112);
CN_in_sigd(2062)	<=	VN_out_sigd(1112);
CN_in_sigd(3062)	<=	VN_out_sigd(1112);
CN_in_sigd(4726)	<=	VN_out_sigd(1112);
CN_in_sigd(894)	<=	VN_out_sigd(1113);
CN_in_sigd(2070)	<=	VN_out_sigd(1113);
CN_in_sigd(3070)	<=	VN_out_sigd(1113);
CN_in_sigd(4734)	<=	VN_out_sigd(1113);
CN_in_sigd(902)	<=	VN_out_sigd(1114);
CN_in_sigd(2078)	<=	VN_out_sigd(1114);
CN_in_sigd(3078)	<=	VN_out_sigd(1114);
CN_in_sigd(4742)	<=	VN_out_sigd(1114);
CN_in_sigd(910)	<=	VN_out_sigd(1115);
CN_in_sigd(2086)	<=	VN_out_sigd(1115);
CN_in_sigd(3086)	<=	VN_out_sigd(1115);
CN_in_sigd(4750)	<=	VN_out_sigd(1115);
CN_in_sigd(918)	<=	VN_out_sigd(1116);
CN_in_sigd(2094)	<=	VN_out_sigd(1116);
CN_in_sigd(3094)	<=	VN_out_sigd(1116);
CN_in_sigd(4326)	<=	VN_out_sigd(1116);
CN_in_sigd(926)	<=	VN_out_sigd(1117);
CN_in_sigd(2102)	<=	VN_out_sigd(1117);
CN_in_sigd(3102)	<=	VN_out_sigd(1117);
CN_in_sigd(4334)	<=	VN_out_sigd(1117);
CN_in_sigd(934)	<=	VN_out_sigd(1118);
CN_in_sigd(2110)	<=	VN_out_sigd(1118);
CN_in_sigd(3110)	<=	VN_out_sigd(1118);
CN_in_sigd(4342)	<=	VN_out_sigd(1118);
CN_in_sigd(942)	<=	VN_out_sigd(1119);
CN_in_sigd(2118)	<=	VN_out_sigd(1119);
CN_in_sigd(3118)	<=	VN_out_sigd(1119);
CN_in_sigd(4350)	<=	VN_out_sigd(1119);
CN_in_sigd(950)	<=	VN_out_sigd(1120);
CN_in_sigd(2126)	<=	VN_out_sigd(1120);
CN_in_sigd(3126)	<=	VN_out_sigd(1120);
CN_in_sigd(4358)	<=	VN_out_sigd(1120);
CN_in_sigd(958)	<=	VN_out_sigd(1121);
CN_in_sigd(2134)	<=	VN_out_sigd(1121);
CN_in_sigd(3134)	<=	VN_out_sigd(1121);
CN_in_sigd(4366)	<=	VN_out_sigd(1121);
CN_in_sigd(966)	<=	VN_out_sigd(1122);
CN_in_sigd(2142)	<=	VN_out_sigd(1122);
CN_in_sigd(3142)	<=	VN_out_sigd(1122);
CN_in_sigd(4374)	<=	VN_out_sigd(1122);
CN_in_sigd(974)	<=	VN_out_sigd(1123);
CN_in_sigd(2150)	<=	VN_out_sigd(1123);
CN_in_sigd(3150)	<=	VN_out_sigd(1123);
CN_in_sigd(4382)	<=	VN_out_sigd(1123);
CN_in_sigd(982)	<=	VN_out_sigd(1124);
CN_in_sigd(2158)	<=	VN_out_sigd(1124);
CN_in_sigd(3158)	<=	VN_out_sigd(1124);
CN_in_sigd(4390)	<=	VN_out_sigd(1124);
CN_in_sigd(990)	<=	VN_out_sigd(1125);
CN_in_sigd(1734)	<=	VN_out_sigd(1125);
CN_in_sigd(3166)	<=	VN_out_sigd(1125);
CN_in_sigd(4398)	<=	VN_out_sigd(1125);
CN_in_sigd(998)	<=	VN_out_sigd(1126);
CN_in_sigd(1742)	<=	VN_out_sigd(1126);
CN_in_sigd(3174)	<=	VN_out_sigd(1126);
CN_in_sigd(4406)	<=	VN_out_sigd(1126);
CN_in_sigd(1006)	<=	VN_out_sigd(1127);
CN_in_sigd(1750)	<=	VN_out_sigd(1127);
CN_in_sigd(3182)	<=	VN_out_sigd(1127);
CN_in_sigd(4414)	<=	VN_out_sigd(1127);
CN_in_sigd(1014)	<=	VN_out_sigd(1128);
CN_in_sigd(1758)	<=	VN_out_sigd(1128);
CN_in_sigd(3190)	<=	VN_out_sigd(1128);
CN_in_sigd(4422)	<=	VN_out_sigd(1128);
CN_in_sigd(1022)	<=	VN_out_sigd(1129);
CN_in_sigd(1766)	<=	VN_out_sigd(1129);
CN_in_sigd(3198)	<=	VN_out_sigd(1129);
CN_in_sigd(4430)	<=	VN_out_sigd(1129);
CN_in_sigd(1030)	<=	VN_out_sigd(1130);
CN_in_sigd(1774)	<=	VN_out_sigd(1130);
CN_in_sigd(3206)	<=	VN_out_sigd(1130);
CN_in_sigd(4438)	<=	VN_out_sigd(1130);
CN_in_sigd(1038)	<=	VN_out_sigd(1131);
CN_in_sigd(1782)	<=	VN_out_sigd(1131);
CN_in_sigd(3214)	<=	VN_out_sigd(1131);
CN_in_sigd(4446)	<=	VN_out_sigd(1131);
CN_in_sigd(1046)	<=	VN_out_sigd(1132);
CN_in_sigd(1790)	<=	VN_out_sigd(1132);
CN_in_sigd(3222)	<=	VN_out_sigd(1132);
CN_in_sigd(4454)	<=	VN_out_sigd(1132);
CN_in_sigd(1054)	<=	VN_out_sigd(1133);
CN_in_sigd(1798)	<=	VN_out_sigd(1133);
CN_in_sigd(3230)	<=	VN_out_sigd(1133);
CN_in_sigd(4462)	<=	VN_out_sigd(1133);
CN_in_sigd(1039)	<=	VN_out_sigd(1134);
CN_in_sigd(2031)	<=	VN_out_sigd(1134);
CN_in_sigd(3135)	<=	VN_out_sigd(1134);
CN_in_sigd(4455)	<=	VN_out_sigd(1134);
CN_in_sigd(1047)	<=	VN_out_sigd(1135);
CN_in_sigd(2039)	<=	VN_out_sigd(1135);
CN_in_sigd(3143)	<=	VN_out_sigd(1135);
CN_in_sigd(4463)	<=	VN_out_sigd(1135);
CN_in_sigd(1055)	<=	VN_out_sigd(1136);
CN_in_sigd(2047)	<=	VN_out_sigd(1136);
CN_in_sigd(3151)	<=	VN_out_sigd(1136);
CN_in_sigd(4471)	<=	VN_out_sigd(1136);
CN_in_sigd(1063)	<=	VN_out_sigd(1137);
CN_in_sigd(2055)	<=	VN_out_sigd(1137);
CN_in_sigd(3159)	<=	VN_out_sigd(1137);
CN_in_sigd(4479)	<=	VN_out_sigd(1137);
CN_in_sigd(1071)	<=	VN_out_sigd(1138);
CN_in_sigd(2063)	<=	VN_out_sigd(1138);
CN_in_sigd(3167)	<=	VN_out_sigd(1138);
CN_in_sigd(4487)	<=	VN_out_sigd(1138);
CN_in_sigd(1079)	<=	VN_out_sigd(1139);
CN_in_sigd(2071)	<=	VN_out_sigd(1139);
CN_in_sigd(3175)	<=	VN_out_sigd(1139);
CN_in_sigd(4495)	<=	VN_out_sigd(1139);
CN_in_sigd(1087)	<=	VN_out_sigd(1140);
CN_in_sigd(2079)	<=	VN_out_sigd(1140);
CN_in_sigd(3183)	<=	VN_out_sigd(1140);
CN_in_sigd(4503)	<=	VN_out_sigd(1140);
CN_in_sigd(1095)	<=	VN_out_sigd(1141);
CN_in_sigd(2087)	<=	VN_out_sigd(1141);
CN_in_sigd(3191)	<=	VN_out_sigd(1141);
CN_in_sigd(4511)	<=	VN_out_sigd(1141);
CN_in_sigd(1103)	<=	VN_out_sigd(1142);
CN_in_sigd(2095)	<=	VN_out_sigd(1142);
CN_in_sigd(3199)	<=	VN_out_sigd(1142);
CN_in_sigd(4519)	<=	VN_out_sigd(1142);
CN_in_sigd(1111)	<=	VN_out_sigd(1143);
CN_in_sigd(2103)	<=	VN_out_sigd(1143);
CN_in_sigd(3207)	<=	VN_out_sigd(1143);
CN_in_sigd(4527)	<=	VN_out_sigd(1143);
CN_in_sigd(1119)	<=	VN_out_sigd(1144);
CN_in_sigd(2111)	<=	VN_out_sigd(1144);
CN_in_sigd(3215)	<=	VN_out_sigd(1144);
CN_in_sigd(4535)	<=	VN_out_sigd(1144);
CN_in_sigd(1127)	<=	VN_out_sigd(1145);
CN_in_sigd(2119)	<=	VN_out_sigd(1145);
CN_in_sigd(3223)	<=	VN_out_sigd(1145);
CN_in_sigd(4543)	<=	VN_out_sigd(1145);
CN_in_sigd(1135)	<=	VN_out_sigd(1146);
CN_in_sigd(2127)	<=	VN_out_sigd(1146);
CN_in_sigd(3231)	<=	VN_out_sigd(1146);
CN_in_sigd(4551)	<=	VN_out_sigd(1146);
CN_in_sigd(1143)	<=	VN_out_sigd(1147);
CN_in_sigd(2135)	<=	VN_out_sigd(1147);
CN_in_sigd(3239)	<=	VN_out_sigd(1147);
CN_in_sigd(4559)	<=	VN_out_sigd(1147);
CN_in_sigd(1151)	<=	VN_out_sigd(1148);
CN_in_sigd(2143)	<=	VN_out_sigd(1148);
CN_in_sigd(3247)	<=	VN_out_sigd(1148);
CN_in_sigd(4567)	<=	VN_out_sigd(1148);
CN_in_sigd(1159)	<=	VN_out_sigd(1149);
CN_in_sigd(2151)	<=	VN_out_sigd(1149);
CN_in_sigd(3255)	<=	VN_out_sigd(1149);
CN_in_sigd(4575)	<=	VN_out_sigd(1149);
CN_in_sigd(1167)	<=	VN_out_sigd(1150);
CN_in_sigd(2159)	<=	VN_out_sigd(1150);
CN_in_sigd(3263)	<=	VN_out_sigd(1150);
CN_in_sigd(4583)	<=	VN_out_sigd(1150);
CN_in_sigd(1175)	<=	VN_out_sigd(1151);
CN_in_sigd(1735)	<=	VN_out_sigd(1151);
CN_in_sigd(3271)	<=	VN_out_sigd(1151);
CN_in_sigd(4591)	<=	VN_out_sigd(1151);
CN_in_sigd(1183)	<=	VN_out_sigd(1152);
CN_in_sigd(1743)	<=	VN_out_sigd(1152);
CN_in_sigd(3279)	<=	VN_out_sigd(1152);
CN_in_sigd(4599)	<=	VN_out_sigd(1152);
CN_in_sigd(1191)	<=	VN_out_sigd(1153);
CN_in_sigd(1751)	<=	VN_out_sigd(1153);
CN_in_sigd(3287)	<=	VN_out_sigd(1153);
CN_in_sigd(4607)	<=	VN_out_sigd(1153);
CN_in_sigd(1199)	<=	VN_out_sigd(1154);
CN_in_sigd(1759)	<=	VN_out_sigd(1154);
CN_in_sigd(3295)	<=	VN_out_sigd(1154);
CN_in_sigd(4615)	<=	VN_out_sigd(1154);
CN_in_sigd(1207)	<=	VN_out_sigd(1155);
CN_in_sigd(1767)	<=	VN_out_sigd(1155);
CN_in_sigd(3303)	<=	VN_out_sigd(1155);
CN_in_sigd(4623)	<=	VN_out_sigd(1155);
CN_in_sigd(1215)	<=	VN_out_sigd(1156);
CN_in_sigd(1775)	<=	VN_out_sigd(1156);
CN_in_sigd(3311)	<=	VN_out_sigd(1156);
CN_in_sigd(4631)	<=	VN_out_sigd(1156);
CN_in_sigd(1223)	<=	VN_out_sigd(1157);
CN_in_sigd(1783)	<=	VN_out_sigd(1157);
CN_in_sigd(3319)	<=	VN_out_sigd(1157);
CN_in_sigd(4639)	<=	VN_out_sigd(1157);
CN_in_sigd(1231)	<=	VN_out_sigd(1158);
CN_in_sigd(1791)	<=	VN_out_sigd(1158);
CN_in_sigd(3327)	<=	VN_out_sigd(1158);
CN_in_sigd(4647)	<=	VN_out_sigd(1158);
CN_in_sigd(1239)	<=	VN_out_sigd(1159);
CN_in_sigd(1799)	<=	VN_out_sigd(1159);
CN_in_sigd(3335)	<=	VN_out_sigd(1159);
CN_in_sigd(4655)	<=	VN_out_sigd(1159);
CN_in_sigd(1247)	<=	VN_out_sigd(1160);
CN_in_sigd(1807)	<=	VN_out_sigd(1160);
CN_in_sigd(3343)	<=	VN_out_sigd(1160);
CN_in_sigd(4663)	<=	VN_out_sigd(1160);
CN_in_sigd(1255)	<=	VN_out_sigd(1161);
CN_in_sigd(1815)	<=	VN_out_sigd(1161);
CN_in_sigd(3351)	<=	VN_out_sigd(1161);
CN_in_sigd(4671)	<=	VN_out_sigd(1161);
CN_in_sigd(1263)	<=	VN_out_sigd(1162);
CN_in_sigd(1823)	<=	VN_out_sigd(1162);
CN_in_sigd(3359)	<=	VN_out_sigd(1162);
CN_in_sigd(4679)	<=	VN_out_sigd(1162);
CN_in_sigd(1271)	<=	VN_out_sigd(1163);
CN_in_sigd(1831)	<=	VN_out_sigd(1163);
CN_in_sigd(3367)	<=	VN_out_sigd(1163);
CN_in_sigd(4687)	<=	VN_out_sigd(1163);
CN_in_sigd(1279)	<=	VN_out_sigd(1164);
CN_in_sigd(1839)	<=	VN_out_sigd(1164);
CN_in_sigd(3375)	<=	VN_out_sigd(1164);
CN_in_sigd(4695)	<=	VN_out_sigd(1164);
CN_in_sigd(1287)	<=	VN_out_sigd(1165);
CN_in_sigd(1847)	<=	VN_out_sigd(1165);
CN_in_sigd(3383)	<=	VN_out_sigd(1165);
CN_in_sigd(4703)	<=	VN_out_sigd(1165);
CN_in_sigd(1295)	<=	VN_out_sigd(1166);
CN_in_sigd(1855)	<=	VN_out_sigd(1166);
CN_in_sigd(3391)	<=	VN_out_sigd(1166);
CN_in_sigd(4711)	<=	VN_out_sigd(1166);
CN_in_sigd(871)	<=	VN_out_sigd(1167);
CN_in_sigd(1863)	<=	VN_out_sigd(1167);
CN_in_sigd(3399)	<=	VN_out_sigd(1167);
CN_in_sigd(4719)	<=	VN_out_sigd(1167);
CN_in_sigd(879)	<=	VN_out_sigd(1168);
CN_in_sigd(1871)	<=	VN_out_sigd(1168);
CN_in_sigd(3407)	<=	VN_out_sigd(1168);
CN_in_sigd(4727)	<=	VN_out_sigd(1168);
CN_in_sigd(887)	<=	VN_out_sigd(1169);
CN_in_sigd(1879)	<=	VN_out_sigd(1169);
CN_in_sigd(3415)	<=	VN_out_sigd(1169);
CN_in_sigd(4735)	<=	VN_out_sigd(1169);
CN_in_sigd(895)	<=	VN_out_sigd(1170);
CN_in_sigd(1887)	<=	VN_out_sigd(1170);
CN_in_sigd(3423)	<=	VN_out_sigd(1170);
CN_in_sigd(4743)	<=	VN_out_sigd(1170);
CN_in_sigd(903)	<=	VN_out_sigd(1171);
CN_in_sigd(1895)	<=	VN_out_sigd(1171);
CN_in_sigd(3431)	<=	VN_out_sigd(1171);
CN_in_sigd(4751)	<=	VN_out_sigd(1171);
CN_in_sigd(911)	<=	VN_out_sigd(1172);
CN_in_sigd(1903)	<=	VN_out_sigd(1172);
CN_in_sigd(3439)	<=	VN_out_sigd(1172);
CN_in_sigd(4327)	<=	VN_out_sigd(1172);
CN_in_sigd(919)	<=	VN_out_sigd(1173);
CN_in_sigd(1911)	<=	VN_out_sigd(1173);
CN_in_sigd(3447)	<=	VN_out_sigd(1173);
CN_in_sigd(4335)	<=	VN_out_sigd(1173);
CN_in_sigd(927)	<=	VN_out_sigd(1174);
CN_in_sigd(1919)	<=	VN_out_sigd(1174);
CN_in_sigd(3455)	<=	VN_out_sigd(1174);
CN_in_sigd(4343)	<=	VN_out_sigd(1174);
CN_in_sigd(935)	<=	VN_out_sigd(1175);
CN_in_sigd(1927)	<=	VN_out_sigd(1175);
CN_in_sigd(3031)	<=	VN_out_sigd(1175);
CN_in_sigd(4351)	<=	VN_out_sigd(1175);
CN_in_sigd(943)	<=	VN_out_sigd(1176);
CN_in_sigd(1935)	<=	VN_out_sigd(1176);
CN_in_sigd(3039)	<=	VN_out_sigd(1176);
CN_in_sigd(4359)	<=	VN_out_sigd(1176);
CN_in_sigd(951)	<=	VN_out_sigd(1177);
CN_in_sigd(1943)	<=	VN_out_sigd(1177);
CN_in_sigd(3047)	<=	VN_out_sigd(1177);
CN_in_sigd(4367)	<=	VN_out_sigd(1177);
CN_in_sigd(959)	<=	VN_out_sigd(1178);
CN_in_sigd(1951)	<=	VN_out_sigd(1178);
CN_in_sigd(3055)	<=	VN_out_sigd(1178);
CN_in_sigd(4375)	<=	VN_out_sigd(1178);
CN_in_sigd(967)	<=	VN_out_sigd(1179);
CN_in_sigd(1959)	<=	VN_out_sigd(1179);
CN_in_sigd(3063)	<=	VN_out_sigd(1179);
CN_in_sigd(4383)	<=	VN_out_sigd(1179);
CN_in_sigd(975)	<=	VN_out_sigd(1180);
CN_in_sigd(1967)	<=	VN_out_sigd(1180);
CN_in_sigd(3071)	<=	VN_out_sigd(1180);
CN_in_sigd(4391)	<=	VN_out_sigd(1180);
CN_in_sigd(983)	<=	VN_out_sigd(1181);
CN_in_sigd(1975)	<=	VN_out_sigd(1181);
CN_in_sigd(3079)	<=	VN_out_sigd(1181);
CN_in_sigd(4399)	<=	VN_out_sigd(1181);
CN_in_sigd(991)	<=	VN_out_sigd(1182);
CN_in_sigd(1983)	<=	VN_out_sigd(1182);
CN_in_sigd(3087)	<=	VN_out_sigd(1182);
CN_in_sigd(4407)	<=	VN_out_sigd(1182);
CN_in_sigd(999)	<=	VN_out_sigd(1183);
CN_in_sigd(1991)	<=	VN_out_sigd(1183);
CN_in_sigd(3095)	<=	VN_out_sigd(1183);
CN_in_sigd(4415)	<=	VN_out_sigd(1183);
CN_in_sigd(1007)	<=	VN_out_sigd(1184);
CN_in_sigd(1999)	<=	VN_out_sigd(1184);
CN_in_sigd(3103)	<=	VN_out_sigd(1184);
CN_in_sigd(4423)	<=	VN_out_sigd(1184);
CN_in_sigd(1015)	<=	VN_out_sigd(1185);
CN_in_sigd(2007)	<=	VN_out_sigd(1185);
CN_in_sigd(3111)	<=	VN_out_sigd(1185);
CN_in_sigd(4431)	<=	VN_out_sigd(1185);
CN_in_sigd(1023)	<=	VN_out_sigd(1186);
CN_in_sigd(2015)	<=	VN_out_sigd(1186);
CN_in_sigd(3119)	<=	VN_out_sigd(1186);
CN_in_sigd(4439)	<=	VN_out_sigd(1186);
CN_in_sigd(1031)	<=	VN_out_sigd(1187);
CN_in_sigd(2023)	<=	VN_out_sigd(1187);
CN_in_sigd(3127)	<=	VN_out_sigd(1187);
CN_in_sigd(4447)	<=	VN_out_sigd(1187);
CN_in_sigd(735)	<=	VN_out_sigd(1188);
CN_in_sigd(2351)	<=	VN_out_sigd(1188);
CN_in_sigd(2719)	<=	VN_out_sigd(1188);
CN_in_sigd(3975)	<=	VN_out_sigd(1188);
CN_in_sigd(743)	<=	VN_out_sigd(1189);
CN_in_sigd(2359)	<=	VN_out_sigd(1189);
CN_in_sigd(2727)	<=	VN_out_sigd(1189);
CN_in_sigd(3983)	<=	VN_out_sigd(1189);
CN_in_sigd(751)	<=	VN_out_sigd(1190);
CN_in_sigd(2367)	<=	VN_out_sigd(1190);
CN_in_sigd(2735)	<=	VN_out_sigd(1190);
CN_in_sigd(3991)	<=	VN_out_sigd(1190);
CN_in_sigd(759)	<=	VN_out_sigd(1191);
CN_in_sigd(2375)	<=	VN_out_sigd(1191);
CN_in_sigd(2743)	<=	VN_out_sigd(1191);
CN_in_sigd(3999)	<=	VN_out_sigd(1191);
CN_in_sigd(767)	<=	VN_out_sigd(1192);
CN_in_sigd(2383)	<=	VN_out_sigd(1192);
CN_in_sigd(2751)	<=	VN_out_sigd(1192);
CN_in_sigd(4007)	<=	VN_out_sigd(1192);
CN_in_sigd(775)	<=	VN_out_sigd(1193);
CN_in_sigd(2391)	<=	VN_out_sigd(1193);
CN_in_sigd(2759)	<=	VN_out_sigd(1193);
CN_in_sigd(4015)	<=	VN_out_sigd(1193);
CN_in_sigd(783)	<=	VN_out_sigd(1194);
CN_in_sigd(2399)	<=	VN_out_sigd(1194);
CN_in_sigd(2767)	<=	VN_out_sigd(1194);
CN_in_sigd(4023)	<=	VN_out_sigd(1194);
CN_in_sigd(791)	<=	VN_out_sigd(1195);
CN_in_sigd(2407)	<=	VN_out_sigd(1195);
CN_in_sigd(2775)	<=	VN_out_sigd(1195);
CN_in_sigd(4031)	<=	VN_out_sigd(1195);
CN_in_sigd(799)	<=	VN_out_sigd(1196);
CN_in_sigd(2415)	<=	VN_out_sigd(1196);
CN_in_sigd(2783)	<=	VN_out_sigd(1196);
CN_in_sigd(4039)	<=	VN_out_sigd(1196);
CN_in_sigd(807)	<=	VN_out_sigd(1197);
CN_in_sigd(2423)	<=	VN_out_sigd(1197);
CN_in_sigd(2791)	<=	VN_out_sigd(1197);
CN_in_sigd(4047)	<=	VN_out_sigd(1197);
CN_in_sigd(815)	<=	VN_out_sigd(1198);
CN_in_sigd(2431)	<=	VN_out_sigd(1198);
CN_in_sigd(2799)	<=	VN_out_sigd(1198);
CN_in_sigd(4055)	<=	VN_out_sigd(1198);
CN_in_sigd(823)	<=	VN_out_sigd(1199);
CN_in_sigd(2439)	<=	VN_out_sigd(1199);
CN_in_sigd(2807)	<=	VN_out_sigd(1199);
CN_in_sigd(4063)	<=	VN_out_sigd(1199);
CN_in_sigd(831)	<=	VN_out_sigd(1200);
CN_in_sigd(2447)	<=	VN_out_sigd(1200);
CN_in_sigd(2815)	<=	VN_out_sigd(1200);
CN_in_sigd(4071)	<=	VN_out_sigd(1200);
CN_in_sigd(839)	<=	VN_out_sigd(1201);
CN_in_sigd(2455)	<=	VN_out_sigd(1201);
CN_in_sigd(2823)	<=	VN_out_sigd(1201);
CN_in_sigd(4079)	<=	VN_out_sigd(1201);
CN_in_sigd(847)	<=	VN_out_sigd(1202);
CN_in_sigd(2463)	<=	VN_out_sigd(1202);
CN_in_sigd(2831)	<=	VN_out_sigd(1202);
CN_in_sigd(4087)	<=	VN_out_sigd(1202);
CN_in_sigd(855)	<=	VN_out_sigd(1203);
CN_in_sigd(2471)	<=	VN_out_sigd(1203);
CN_in_sigd(2839)	<=	VN_out_sigd(1203);
CN_in_sigd(4095)	<=	VN_out_sigd(1203);
CN_in_sigd(863)	<=	VN_out_sigd(1204);
CN_in_sigd(2479)	<=	VN_out_sigd(1204);
CN_in_sigd(2847)	<=	VN_out_sigd(1204);
CN_in_sigd(4103)	<=	VN_out_sigd(1204);
CN_in_sigd(439)	<=	VN_out_sigd(1205);
CN_in_sigd(2487)	<=	VN_out_sigd(1205);
CN_in_sigd(2855)	<=	VN_out_sigd(1205);
CN_in_sigd(4111)	<=	VN_out_sigd(1205);
CN_in_sigd(447)	<=	VN_out_sigd(1206);
CN_in_sigd(2495)	<=	VN_out_sigd(1206);
CN_in_sigd(2863)	<=	VN_out_sigd(1206);
CN_in_sigd(4119)	<=	VN_out_sigd(1206);
CN_in_sigd(455)	<=	VN_out_sigd(1207);
CN_in_sigd(2503)	<=	VN_out_sigd(1207);
CN_in_sigd(2871)	<=	VN_out_sigd(1207);
CN_in_sigd(4127)	<=	VN_out_sigd(1207);
CN_in_sigd(463)	<=	VN_out_sigd(1208);
CN_in_sigd(2511)	<=	VN_out_sigd(1208);
CN_in_sigd(2879)	<=	VN_out_sigd(1208);
CN_in_sigd(4135)	<=	VN_out_sigd(1208);
CN_in_sigd(471)	<=	VN_out_sigd(1209);
CN_in_sigd(2519)	<=	VN_out_sigd(1209);
CN_in_sigd(2887)	<=	VN_out_sigd(1209);
CN_in_sigd(4143)	<=	VN_out_sigd(1209);
CN_in_sigd(479)	<=	VN_out_sigd(1210);
CN_in_sigd(2527)	<=	VN_out_sigd(1210);
CN_in_sigd(2895)	<=	VN_out_sigd(1210);
CN_in_sigd(4151)	<=	VN_out_sigd(1210);
CN_in_sigd(487)	<=	VN_out_sigd(1211);
CN_in_sigd(2535)	<=	VN_out_sigd(1211);
CN_in_sigd(2903)	<=	VN_out_sigd(1211);
CN_in_sigd(4159)	<=	VN_out_sigd(1211);
CN_in_sigd(495)	<=	VN_out_sigd(1212);
CN_in_sigd(2543)	<=	VN_out_sigd(1212);
CN_in_sigd(2911)	<=	VN_out_sigd(1212);
CN_in_sigd(4167)	<=	VN_out_sigd(1212);
CN_in_sigd(503)	<=	VN_out_sigd(1213);
CN_in_sigd(2551)	<=	VN_out_sigd(1213);
CN_in_sigd(2919)	<=	VN_out_sigd(1213);
CN_in_sigd(4175)	<=	VN_out_sigd(1213);
CN_in_sigd(511)	<=	VN_out_sigd(1214);
CN_in_sigd(2559)	<=	VN_out_sigd(1214);
CN_in_sigd(2927)	<=	VN_out_sigd(1214);
CN_in_sigd(4183)	<=	VN_out_sigd(1214);
CN_in_sigd(519)	<=	VN_out_sigd(1215);
CN_in_sigd(2567)	<=	VN_out_sigd(1215);
CN_in_sigd(2935)	<=	VN_out_sigd(1215);
CN_in_sigd(4191)	<=	VN_out_sigd(1215);
CN_in_sigd(527)	<=	VN_out_sigd(1216);
CN_in_sigd(2575)	<=	VN_out_sigd(1216);
CN_in_sigd(2943)	<=	VN_out_sigd(1216);
CN_in_sigd(4199)	<=	VN_out_sigd(1216);
CN_in_sigd(535)	<=	VN_out_sigd(1217);
CN_in_sigd(2583)	<=	VN_out_sigd(1217);
CN_in_sigd(2951)	<=	VN_out_sigd(1217);
CN_in_sigd(4207)	<=	VN_out_sigd(1217);
CN_in_sigd(543)	<=	VN_out_sigd(1218);
CN_in_sigd(2591)	<=	VN_out_sigd(1218);
CN_in_sigd(2959)	<=	VN_out_sigd(1218);
CN_in_sigd(4215)	<=	VN_out_sigd(1218);
CN_in_sigd(551)	<=	VN_out_sigd(1219);
CN_in_sigd(2167)	<=	VN_out_sigd(1219);
CN_in_sigd(2967)	<=	VN_out_sigd(1219);
CN_in_sigd(4223)	<=	VN_out_sigd(1219);
CN_in_sigd(559)	<=	VN_out_sigd(1220);
CN_in_sigd(2175)	<=	VN_out_sigd(1220);
CN_in_sigd(2975)	<=	VN_out_sigd(1220);
CN_in_sigd(4231)	<=	VN_out_sigd(1220);
CN_in_sigd(567)	<=	VN_out_sigd(1221);
CN_in_sigd(2183)	<=	VN_out_sigd(1221);
CN_in_sigd(2983)	<=	VN_out_sigd(1221);
CN_in_sigd(4239)	<=	VN_out_sigd(1221);
CN_in_sigd(575)	<=	VN_out_sigd(1222);
CN_in_sigd(2191)	<=	VN_out_sigd(1222);
CN_in_sigd(2991)	<=	VN_out_sigd(1222);
CN_in_sigd(4247)	<=	VN_out_sigd(1222);
CN_in_sigd(583)	<=	VN_out_sigd(1223);
CN_in_sigd(2199)	<=	VN_out_sigd(1223);
CN_in_sigd(2999)	<=	VN_out_sigd(1223);
CN_in_sigd(4255)	<=	VN_out_sigd(1223);
CN_in_sigd(591)	<=	VN_out_sigd(1224);
CN_in_sigd(2207)	<=	VN_out_sigd(1224);
CN_in_sigd(3007)	<=	VN_out_sigd(1224);
CN_in_sigd(4263)	<=	VN_out_sigd(1224);
CN_in_sigd(599)	<=	VN_out_sigd(1225);
CN_in_sigd(2215)	<=	VN_out_sigd(1225);
CN_in_sigd(3015)	<=	VN_out_sigd(1225);
CN_in_sigd(4271)	<=	VN_out_sigd(1225);
CN_in_sigd(607)	<=	VN_out_sigd(1226);
CN_in_sigd(2223)	<=	VN_out_sigd(1226);
CN_in_sigd(3023)	<=	VN_out_sigd(1226);
CN_in_sigd(4279)	<=	VN_out_sigd(1226);
CN_in_sigd(615)	<=	VN_out_sigd(1227);
CN_in_sigd(2231)	<=	VN_out_sigd(1227);
CN_in_sigd(2599)	<=	VN_out_sigd(1227);
CN_in_sigd(4287)	<=	VN_out_sigd(1227);
CN_in_sigd(623)	<=	VN_out_sigd(1228);
CN_in_sigd(2239)	<=	VN_out_sigd(1228);
CN_in_sigd(2607)	<=	VN_out_sigd(1228);
CN_in_sigd(4295)	<=	VN_out_sigd(1228);
CN_in_sigd(631)	<=	VN_out_sigd(1229);
CN_in_sigd(2247)	<=	VN_out_sigd(1229);
CN_in_sigd(2615)	<=	VN_out_sigd(1229);
CN_in_sigd(4303)	<=	VN_out_sigd(1229);
CN_in_sigd(639)	<=	VN_out_sigd(1230);
CN_in_sigd(2255)	<=	VN_out_sigd(1230);
CN_in_sigd(2623)	<=	VN_out_sigd(1230);
CN_in_sigd(4311)	<=	VN_out_sigd(1230);
CN_in_sigd(647)	<=	VN_out_sigd(1231);
CN_in_sigd(2263)	<=	VN_out_sigd(1231);
CN_in_sigd(2631)	<=	VN_out_sigd(1231);
CN_in_sigd(4319)	<=	VN_out_sigd(1231);
CN_in_sigd(655)	<=	VN_out_sigd(1232);
CN_in_sigd(2271)	<=	VN_out_sigd(1232);
CN_in_sigd(2639)	<=	VN_out_sigd(1232);
CN_in_sigd(3895)	<=	VN_out_sigd(1232);
CN_in_sigd(663)	<=	VN_out_sigd(1233);
CN_in_sigd(2279)	<=	VN_out_sigd(1233);
CN_in_sigd(2647)	<=	VN_out_sigd(1233);
CN_in_sigd(3903)	<=	VN_out_sigd(1233);
CN_in_sigd(671)	<=	VN_out_sigd(1234);
CN_in_sigd(2287)	<=	VN_out_sigd(1234);
CN_in_sigd(2655)	<=	VN_out_sigd(1234);
CN_in_sigd(3911)	<=	VN_out_sigd(1234);
CN_in_sigd(679)	<=	VN_out_sigd(1235);
CN_in_sigd(2295)	<=	VN_out_sigd(1235);
CN_in_sigd(2663)	<=	VN_out_sigd(1235);
CN_in_sigd(3919)	<=	VN_out_sigd(1235);
CN_in_sigd(687)	<=	VN_out_sigd(1236);
CN_in_sigd(2303)	<=	VN_out_sigd(1236);
CN_in_sigd(2671)	<=	VN_out_sigd(1236);
CN_in_sigd(3927)	<=	VN_out_sigd(1236);
CN_in_sigd(695)	<=	VN_out_sigd(1237);
CN_in_sigd(2311)	<=	VN_out_sigd(1237);
CN_in_sigd(2679)	<=	VN_out_sigd(1237);
CN_in_sigd(3935)	<=	VN_out_sigd(1237);
CN_in_sigd(703)	<=	VN_out_sigd(1238);
CN_in_sigd(2319)	<=	VN_out_sigd(1238);
CN_in_sigd(2687)	<=	VN_out_sigd(1238);
CN_in_sigd(3943)	<=	VN_out_sigd(1238);
CN_in_sigd(711)	<=	VN_out_sigd(1239);
CN_in_sigd(2327)	<=	VN_out_sigd(1239);
CN_in_sigd(2695)	<=	VN_out_sigd(1239);
CN_in_sigd(3951)	<=	VN_out_sigd(1239);
CN_in_sigd(719)	<=	VN_out_sigd(1240);
CN_in_sigd(2335)	<=	VN_out_sigd(1240);
CN_in_sigd(2703)	<=	VN_out_sigd(1240);
CN_in_sigd(3959)	<=	VN_out_sigd(1240);
CN_in_sigd(727)	<=	VN_out_sigd(1241);
CN_in_sigd(2343)	<=	VN_out_sigd(1241);
CN_in_sigd(2711)	<=	VN_out_sigd(1241);
CN_in_sigd(3967)	<=	VN_out_sigd(1241);
CN_in_sigd(7)	<=	VN_out_sigd(1242);
CN_in_sigd(1519)	<=	VN_out_sigd(1242);
CN_in_sigd(3567)	<=	VN_out_sigd(1242);
CN_in_sigd(5071)	<=	VN_out_sigd(1242);
CN_in_sigd(15)	<=	VN_out_sigd(1243);
CN_in_sigd(1527)	<=	VN_out_sigd(1243);
CN_in_sigd(3575)	<=	VN_out_sigd(1243);
CN_in_sigd(5079)	<=	VN_out_sigd(1243);
CN_in_sigd(23)	<=	VN_out_sigd(1244);
CN_in_sigd(1535)	<=	VN_out_sigd(1244);
CN_in_sigd(3583)	<=	VN_out_sigd(1244);
CN_in_sigd(5087)	<=	VN_out_sigd(1244);
CN_in_sigd(31)	<=	VN_out_sigd(1245);
CN_in_sigd(1543)	<=	VN_out_sigd(1245);
CN_in_sigd(3591)	<=	VN_out_sigd(1245);
CN_in_sigd(5095)	<=	VN_out_sigd(1245);
CN_in_sigd(39)	<=	VN_out_sigd(1246);
CN_in_sigd(1551)	<=	VN_out_sigd(1246);
CN_in_sigd(3599)	<=	VN_out_sigd(1246);
CN_in_sigd(5103)	<=	VN_out_sigd(1246);
CN_in_sigd(47)	<=	VN_out_sigd(1247);
CN_in_sigd(1559)	<=	VN_out_sigd(1247);
CN_in_sigd(3607)	<=	VN_out_sigd(1247);
CN_in_sigd(5111)	<=	VN_out_sigd(1247);
CN_in_sigd(55)	<=	VN_out_sigd(1248);
CN_in_sigd(1567)	<=	VN_out_sigd(1248);
CN_in_sigd(3615)	<=	VN_out_sigd(1248);
CN_in_sigd(5119)	<=	VN_out_sigd(1248);
CN_in_sigd(63)	<=	VN_out_sigd(1249);
CN_in_sigd(1575)	<=	VN_out_sigd(1249);
CN_in_sigd(3623)	<=	VN_out_sigd(1249);
CN_in_sigd(5127)	<=	VN_out_sigd(1249);
CN_in_sigd(71)	<=	VN_out_sigd(1250);
CN_in_sigd(1583)	<=	VN_out_sigd(1250);
CN_in_sigd(3631)	<=	VN_out_sigd(1250);
CN_in_sigd(5135)	<=	VN_out_sigd(1250);
CN_in_sigd(79)	<=	VN_out_sigd(1251);
CN_in_sigd(1591)	<=	VN_out_sigd(1251);
CN_in_sigd(3639)	<=	VN_out_sigd(1251);
CN_in_sigd(5143)	<=	VN_out_sigd(1251);
CN_in_sigd(87)	<=	VN_out_sigd(1252);
CN_in_sigd(1599)	<=	VN_out_sigd(1252);
CN_in_sigd(3647)	<=	VN_out_sigd(1252);
CN_in_sigd(5151)	<=	VN_out_sigd(1252);
CN_in_sigd(95)	<=	VN_out_sigd(1253);
CN_in_sigd(1607)	<=	VN_out_sigd(1253);
CN_in_sigd(3655)	<=	VN_out_sigd(1253);
CN_in_sigd(5159)	<=	VN_out_sigd(1253);
CN_in_sigd(103)	<=	VN_out_sigd(1254);
CN_in_sigd(1615)	<=	VN_out_sigd(1254);
CN_in_sigd(3663)	<=	VN_out_sigd(1254);
CN_in_sigd(5167)	<=	VN_out_sigd(1254);
CN_in_sigd(111)	<=	VN_out_sigd(1255);
CN_in_sigd(1623)	<=	VN_out_sigd(1255);
CN_in_sigd(3671)	<=	VN_out_sigd(1255);
CN_in_sigd(5175)	<=	VN_out_sigd(1255);
CN_in_sigd(119)	<=	VN_out_sigd(1256);
CN_in_sigd(1631)	<=	VN_out_sigd(1256);
CN_in_sigd(3679)	<=	VN_out_sigd(1256);
CN_in_sigd(5183)	<=	VN_out_sigd(1256);
CN_in_sigd(127)	<=	VN_out_sigd(1257);
CN_in_sigd(1639)	<=	VN_out_sigd(1257);
CN_in_sigd(3687)	<=	VN_out_sigd(1257);
CN_in_sigd(4759)	<=	VN_out_sigd(1257);
CN_in_sigd(135)	<=	VN_out_sigd(1258);
CN_in_sigd(1647)	<=	VN_out_sigd(1258);
CN_in_sigd(3695)	<=	VN_out_sigd(1258);
CN_in_sigd(4767)	<=	VN_out_sigd(1258);
CN_in_sigd(143)	<=	VN_out_sigd(1259);
CN_in_sigd(1655)	<=	VN_out_sigd(1259);
CN_in_sigd(3703)	<=	VN_out_sigd(1259);
CN_in_sigd(4775)	<=	VN_out_sigd(1259);
CN_in_sigd(151)	<=	VN_out_sigd(1260);
CN_in_sigd(1663)	<=	VN_out_sigd(1260);
CN_in_sigd(3711)	<=	VN_out_sigd(1260);
CN_in_sigd(4783)	<=	VN_out_sigd(1260);
CN_in_sigd(159)	<=	VN_out_sigd(1261);
CN_in_sigd(1671)	<=	VN_out_sigd(1261);
CN_in_sigd(3719)	<=	VN_out_sigd(1261);
CN_in_sigd(4791)	<=	VN_out_sigd(1261);
CN_in_sigd(167)	<=	VN_out_sigd(1262);
CN_in_sigd(1679)	<=	VN_out_sigd(1262);
CN_in_sigd(3727)	<=	VN_out_sigd(1262);
CN_in_sigd(4799)	<=	VN_out_sigd(1262);
CN_in_sigd(175)	<=	VN_out_sigd(1263);
CN_in_sigd(1687)	<=	VN_out_sigd(1263);
CN_in_sigd(3735)	<=	VN_out_sigd(1263);
CN_in_sigd(4807)	<=	VN_out_sigd(1263);
CN_in_sigd(183)	<=	VN_out_sigd(1264);
CN_in_sigd(1695)	<=	VN_out_sigd(1264);
CN_in_sigd(3743)	<=	VN_out_sigd(1264);
CN_in_sigd(4815)	<=	VN_out_sigd(1264);
CN_in_sigd(191)	<=	VN_out_sigd(1265);
CN_in_sigd(1703)	<=	VN_out_sigd(1265);
CN_in_sigd(3751)	<=	VN_out_sigd(1265);
CN_in_sigd(4823)	<=	VN_out_sigd(1265);
CN_in_sigd(199)	<=	VN_out_sigd(1266);
CN_in_sigd(1711)	<=	VN_out_sigd(1266);
CN_in_sigd(3759)	<=	VN_out_sigd(1266);
CN_in_sigd(4831)	<=	VN_out_sigd(1266);
CN_in_sigd(207)	<=	VN_out_sigd(1267);
CN_in_sigd(1719)	<=	VN_out_sigd(1267);
CN_in_sigd(3767)	<=	VN_out_sigd(1267);
CN_in_sigd(4839)	<=	VN_out_sigd(1267);
CN_in_sigd(215)	<=	VN_out_sigd(1268);
CN_in_sigd(1727)	<=	VN_out_sigd(1268);
CN_in_sigd(3775)	<=	VN_out_sigd(1268);
CN_in_sigd(4847)	<=	VN_out_sigd(1268);
CN_in_sigd(223)	<=	VN_out_sigd(1269);
CN_in_sigd(1303)	<=	VN_out_sigd(1269);
CN_in_sigd(3783)	<=	VN_out_sigd(1269);
CN_in_sigd(4855)	<=	VN_out_sigd(1269);
CN_in_sigd(231)	<=	VN_out_sigd(1270);
CN_in_sigd(1311)	<=	VN_out_sigd(1270);
CN_in_sigd(3791)	<=	VN_out_sigd(1270);
CN_in_sigd(4863)	<=	VN_out_sigd(1270);
CN_in_sigd(239)	<=	VN_out_sigd(1271);
CN_in_sigd(1319)	<=	VN_out_sigd(1271);
CN_in_sigd(3799)	<=	VN_out_sigd(1271);
CN_in_sigd(4871)	<=	VN_out_sigd(1271);
CN_in_sigd(247)	<=	VN_out_sigd(1272);
CN_in_sigd(1327)	<=	VN_out_sigd(1272);
CN_in_sigd(3807)	<=	VN_out_sigd(1272);
CN_in_sigd(4879)	<=	VN_out_sigd(1272);
CN_in_sigd(255)	<=	VN_out_sigd(1273);
CN_in_sigd(1335)	<=	VN_out_sigd(1273);
CN_in_sigd(3815)	<=	VN_out_sigd(1273);
CN_in_sigd(4887)	<=	VN_out_sigd(1273);
CN_in_sigd(263)	<=	VN_out_sigd(1274);
CN_in_sigd(1343)	<=	VN_out_sigd(1274);
CN_in_sigd(3823)	<=	VN_out_sigd(1274);
CN_in_sigd(4895)	<=	VN_out_sigd(1274);
CN_in_sigd(271)	<=	VN_out_sigd(1275);
CN_in_sigd(1351)	<=	VN_out_sigd(1275);
CN_in_sigd(3831)	<=	VN_out_sigd(1275);
CN_in_sigd(4903)	<=	VN_out_sigd(1275);
CN_in_sigd(279)	<=	VN_out_sigd(1276);
CN_in_sigd(1359)	<=	VN_out_sigd(1276);
CN_in_sigd(3839)	<=	VN_out_sigd(1276);
CN_in_sigd(4911)	<=	VN_out_sigd(1276);
CN_in_sigd(287)	<=	VN_out_sigd(1277);
CN_in_sigd(1367)	<=	VN_out_sigd(1277);
CN_in_sigd(3847)	<=	VN_out_sigd(1277);
CN_in_sigd(4919)	<=	VN_out_sigd(1277);
CN_in_sigd(295)	<=	VN_out_sigd(1278);
CN_in_sigd(1375)	<=	VN_out_sigd(1278);
CN_in_sigd(3855)	<=	VN_out_sigd(1278);
CN_in_sigd(4927)	<=	VN_out_sigd(1278);
CN_in_sigd(303)	<=	VN_out_sigd(1279);
CN_in_sigd(1383)	<=	VN_out_sigd(1279);
CN_in_sigd(3863)	<=	VN_out_sigd(1279);
CN_in_sigd(4935)	<=	VN_out_sigd(1279);
CN_in_sigd(311)	<=	VN_out_sigd(1280);
CN_in_sigd(1391)	<=	VN_out_sigd(1280);
CN_in_sigd(3871)	<=	VN_out_sigd(1280);
CN_in_sigd(4943)	<=	VN_out_sigd(1280);
CN_in_sigd(319)	<=	VN_out_sigd(1281);
CN_in_sigd(1399)	<=	VN_out_sigd(1281);
CN_in_sigd(3879)	<=	VN_out_sigd(1281);
CN_in_sigd(4951)	<=	VN_out_sigd(1281);
CN_in_sigd(327)	<=	VN_out_sigd(1282);
CN_in_sigd(1407)	<=	VN_out_sigd(1282);
CN_in_sigd(3887)	<=	VN_out_sigd(1282);
CN_in_sigd(4959)	<=	VN_out_sigd(1282);
CN_in_sigd(335)	<=	VN_out_sigd(1283);
CN_in_sigd(1415)	<=	VN_out_sigd(1283);
CN_in_sigd(3463)	<=	VN_out_sigd(1283);
CN_in_sigd(4967)	<=	VN_out_sigd(1283);
CN_in_sigd(343)	<=	VN_out_sigd(1284);
CN_in_sigd(1423)	<=	VN_out_sigd(1284);
CN_in_sigd(3471)	<=	VN_out_sigd(1284);
CN_in_sigd(4975)	<=	VN_out_sigd(1284);
CN_in_sigd(351)	<=	VN_out_sigd(1285);
CN_in_sigd(1431)	<=	VN_out_sigd(1285);
CN_in_sigd(3479)	<=	VN_out_sigd(1285);
CN_in_sigd(4983)	<=	VN_out_sigd(1285);
CN_in_sigd(359)	<=	VN_out_sigd(1286);
CN_in_sigd(1439)	<=	VN_out_sigd(1286);
CN_in_sigd(3487)	<=	VN_out_sigd(1286);
CN_in_sigd(4991)	<=	VN_out_sigd(1286);
CN_in_sigd(367)	<=	VN_out_sigd(1287);
CN_in_sigd(1447)	<=	VN_out_sigd(1287);
CN_in_sigd(3495)	<=	VN_out_sigd(1287);
CN_in_sigd(4999)	<=	VN_out_sigd(1287);
CN_in_sigd(375)	<=	VN_out_sigd(1288);
CN_in_sigd(1455)	<=	VN_out_sigd(1288);
CN_in_sigd(3503)	<=	VN_out_sigd(1288);
CN_in_sigd(5007)	<=	VN_out_sigd(1288);
CN_in_sigd(383)	<=	VN_out_sigd(1289);
CN_in_sigd(1463)	<=	VN_out_sigd(1289);
CN_in_sigd(3511)	<=	VN_out_sigd(1289);
CN_in_sigd(5015)	<=	VN_out_sigd(1289);
CN_in_sigd(391)	<=	VN_out_sigd(1290);
CN_in_sigd(1471)	<=	VN_out_sigd(1290);
CN_in_sigd(3519)	<=	VN_out_sigd(1290);
CN_in_sigd(5023)	<=	VN_out_sigd(1290);
CN_in_sigd(399)	<=	VN_out_sigd(1291);
CN_in_sigd(1479)	<=	VN_out_sigd(1291);
CN_in_sigd(3527)	<=	VN_out_sigd(1291);
CN_in_sigd(5031)	<=	VN_out_sigd(1291);
CN_in_sigd(407)	<=	VN_out_sigd(1292);
CN_in_sigd(1487)	<=	VN_out_sigd(1292);
CN_in_sigd(3535)	<=	VN_out_sigd(1292);
CN_in_sigd(5039)	<=	VN_out_sigd(1292);
CN_in_sigd(415)	<=	VN_out_sigd(1293);
CN_in_sigd(1495)	<=	VN_out_sigd(1293);
CN_in_sigd(3543)	<=	VN_out_sigd(1293);
CN_in_sigd(5047)	<=	VN_out_sigd(1293);
CN_in_sigd(423)	<=	VN_out_sigd(1294);
CN_in_sigd(1503)	<=	VN_out_sigd(1294);
CN_in_sigd(3551)	<=	VN_out_sigd(1294);
CN_in_sigd(5055)	<=	VN_out_sigd(1294);
CN_in_sigd(431)	<=	VN_out_sigd(1295);
CN_in_sigd(1511)	<=	VN_out_sigd(1295);
CN_in_sigd(3559)	<=	VN_out_sigd(1295);
CN_in_sigd(5063)	<=	VN_out_sigd(1295);



VN_in_sig(44)	<=	CN_out_sig(0);
VN_in_sig(972)	<=	CN_out_sig(1);
VN_in_sig(1860)	<=	CN_out_sig(2);
VN_in_sig(2008)	<=	CN_out_sig(3);
VN_in_sig(2984)	<=	CN_out_sig(4);
VN_in_sig(3632)	<=	CN_out_sig(5);
VN_in_sig(3920)	<=	CN_out_sig(6);
VN_in_sig(4968)	<=	CN_out_sig(7);
VN_in_sig(48)	<=	CN_out_sig(8);
VN_in_sig(976)	<=	CN_out_sig(9);
VN_in_sig(1864)	<=	CN_out_sig(10);
VN_in_sig(2012)	<=	CN_out_sig(11);
VN_in_sig(2988)	<=	CN_out_sig(12);
VN_in_sig(3636)	<=	CN_out_sig(13);
VN_in_sig(3924)	<=	CN_out_sig(14);
VN_in_sig(4972)	<=	CN_out_sig(15);
VN_in_sig(52)	<=	CN_out_sig(16);
VN_in_sig(980)	<=	CN_out_sig(17);
VN_in_sig(1868)	<=	CN_out_sig(18);
VN_in_sig(2016)	<=	CN_out_sig(19);
VN_in_sig(2992)	<=	CN_out_sig(20);
VN_in_sig(3640)	<=	CN_out_sig(21);
VN_in_sig(3928)	<=	CN_out_sig(22);
VN_in_sig(4976)	<=	CN_out_sig(23);
VN_in_sig(56)	<=	CN_out_sig(24);
VN_in_sig(984)	<=	CN_out_sig(25);
VN_in_sig(1872)	<=	CN_out_sig(26);
VN_in_sig(2020)	<=	CN_out_sig(27);
VN_in_sig(2996)	<=	CN_out_sig(28);
VN_in_sig(3644)	<=	CN_out_sig(29);
VN_in_sig(3932)	<=	CN_out_sig(30);
VN_in_sig(4980)	<=	CN_out_sig(31);
VN_in_sig(60)	<=	CN_out_sig(32);
VN_in_sig(988)	<=	CN_out_sig(33);
VN_in_sig(1876)	<=	CN_out_sig(34);
VN_in_sig(2024)	<=	CN_out_sig(35);
VN_in_sig(3000)	<=	CN_out_sig(36);
VN_in_sig(3648)	<=	CN_out_sig(37);
VN_in_sig(3936)	<=	CN_out_sig(38);
VN_in_sig(4984)	<=	CN_out_sig(39);
VN_in_sig(64)	<=	CN_out_sig(40);
VN_in_sig(992)	<=	CN_out_sig(41);
VN_in_sig(1880)	<=	CN_out_sig(42);
VN_in_sig(2028)	<=	CN_out_sig(43);
VN_in_sig(3004)	<=	CN_out_sig(44);
VN_in_sig(3652)	<=	CN_out_sig(45);
VN_in_sig(3940)	<=	CN_out_sig(46);
VN_in_sig(4988)	<=	CN_out_sig(47);
VN_in_sig(68)	<=	CN_out_sig(48);
VN_in_sig(996)	<=	CN_out_sig(49);
VN_in_sig(1884)	<=	CN_out_sig(50);
VN_in_sig(2032)	<=	CN_out_sig(51);
VN_in_sig(3008)	<=	CN_out_sig(52);
VN_in_sig(3656)	<=	CN_out_sig(53);
VN_in_sig(3944)	<=	CN_out_sig(54);
VN_in_sig(4992)	<=	CN_out_sig(55);
VN_in_sig(72)	<=	CN_out_sig(56);
VN_in_sig(1000)	<=	CN_out_sig(57);
VN_in_sig(1888)	<=	CN_out_sig(58);
VN_in_sig(2036)	<=	CN_out_sig(59);
VN_in_sig(3012)	<=	CN_out_sig(60);
VN_in_sig(3660)	<=	CN_out_sig(61);
VN_in_sig(3948)	<=	CN_out_sig(62);
VN_in_sig(4996)	<=	CN_out_sig(63);
VN_in_sig(76)	<=	CN_out_sig(64);
VN_in_sig(1004)	<=	CN_out_sig(65);
VN_in_sig(1892)	<=	CN_out_sig(66);
VN_in_sig(2040)	<=	CN_out_sig(67);
VN_in_sig(3016)	<=	CN_out_sig(68);
VN_in_sig(3664)	<=	CN_out_sig(69);
VN_in_sig(3952)	<=	CN_out_sig(70);
VN_in_sig(5000)	<=	CN_out_sig(71);
VN_in_sig(80)	<=	CN_out_sig(72);
VN_in_sig(1008)	<=	CN_out_sig(73);
VN_in_sig(1896)	<=	CN_out_sig(74);
VN_in_sig(2044)	<=	CN_out_sig(75);
VN_in_sig(3020)	<=	CN_out_sig(76);
VN_in_sig(3668)	<=	CN_out_sig(77);
VN_in_sig(3956)	<=	CN_out_sig(78);
VN_in_sig(5004)	<=	CN_out_sig(79);
VN_in_sig(84)	<=	CN_out_sig(80);
VN_in_sig(1012)	<=	CN_out_sig(81);
VN_in_sig(1900)	<=	CN_out_sig(82);
VN_in_sig(2048)	<=	CN_out_sig(83);
VN_in_sig(2808)	<=	CN_out_sig(84);
VN_in_sig(3456)	<=	CN_out_sig(85);
VN_in_sig(3960)	<=	CN_out_sig(86);
VN_in_sig(5008)	<=	CN_out_sig(87);
VN_in_sig(88)	<=	CN_out_sig(88);
VN_in_sig(1016)	<=	CN_out_sig(89);
VN_in_sig(1904)	<=	CN_out_sig(90);
VN_in_sig(2052)	<=	CN_out_sig(91);
VN_in_sig(2812)	<=	CN_out_sig(92);
VN_in_sig(3460)	<=	CN_out_sig(93);
VN_in_sig(3964)	<=	CN_out_sig(94);
VN_in_sig(5012)	<=	CN_out_sig(95);
VN_in_sig(92)	<=	CN_out_sig(96);
VN_in_sig(1020)	<=	CN_out_sig(97);
VN_in_sig(1908)	<=	CN_out_sig(98);
VN_in_sig(2056)	<=	CN_out_sig(99);
VN_in_sig(2816)	<=	CN_out_sig(100);
VN_in_sig(3464)	<=	CN_out_sig(101);
VN_in_sig(3968)	<=	CN_out_sig(102);
VN_in_sig(5016)	<=	CN_out_sig(103);
VN_in_sig(96)	<=	CN_out_sig(104);
VN_in_sig(1024)	<=	CN_out_sig(105);
VN_in_sig(1912)	<=	CN_out_sig(106);
VN_in_sig(2060)	<=	CN_out_sig(107);
VN_in_sig(2820)	<=	CN_out_sig(108);
VN_in_sig(3468)	<=	CN_out_sig(109);
VN_in_sig(3972)	<=	CN_out_sig(110);
VN_in_sig(5020)	<=	CN_out_sig(111);
VN_in_sig(100)	<=	CN_out_sig(112);
VN_in_sig(1028)	<=	CN_out_sig(113);
VN_in_sig(1916)	<=	CN_out_sig(114);
VN_in_sig(2064)	<=	CN_out_sig(115);
VN_in_sig(2824)	<=	CN_out_sig(116);
VN_in_sig(3472)	<=	CN_out_sig(117);
VN_in_sig(3976)	<=	CN_out_sig(118);
VN_in_sig(5024)	<=	CN_out_sig(119);
VN_in_sig(104)	<=	CN_out_sig(120);
VN_in_sig(1032)	<=	CN_out_sig(121);
VN_in_sig(1920)	<=	CN_out_sig(122);
VN_in_sig(2068)	<=	CN_out_sig(123);
VN_in_sig(2828)	<=	CN_out_sig(124);
VN_in_sig(3476)	<=	CN_out_sig(125);
VN_in_sig(3980)	<=	CN_out_sig(126);
VN_in_sig(5028)	<=	CN_out_sig(127);
VN_in_sig(108)	<=	CN_out_sig(128);
VN_in_sig(1036)	<=	CN_out_sig(129);
VN_in_sig(1924)	<=	CN_out_sig(130);
VN_in_sig(2072)	<=	CN_out_sig(131);
VN_in_sig(2832)	<=	CN_out_sig(132);
VN_in_sig(3480)	<=	CN_out_sig(133);
VN_in_sig(3984)	<=	CN_out_sig(134);
VN_in_sig(5032)	<=	CN_out_sig(135);
VN_in_sig(112)	<=	CN_out_sig(136);
VN_in_sig(1040)	<=	CN_out_sig(137);
VN_in_sig(1928)	<=	CN_out_sig(138);
VN_in_sig(2076)	<=	CN_out_sig(139);
VN_in_sig(2836)	<=	CN_out_sig(140);
VN_in_sig(3484)	<=	CN_out_sig(141);
VN_in_sig(3988)	<=	CN_out_sig(142);
VN_in_sig(5036)	<=	CN_out_sig(143);
VN_in_sig(116)	<=	CN_out_sig(144);
VN_in_sig(1044)	<=	CN_out_sig(145);
VN_in_sig(1932)	<=	CN_out_sig(146);
VN_in_sig(2080)	<=	CN_out_sig(147);
VN_in_sig(2840)	<=	CN_out_sig(148);
VN_in_sig(3488)	<=	CN_out_sig(149);
VN_in_sig(3992)	<=	CN_out_sig(150);
VN_in_sig(5040)	<=	CN_out_sig(151);
VN_in_sig(120)	<=	CN_out_sig(152);
VN_in_sig(1048)	<=	CN_out_sig(153);
VN_in_sig(1936)	<=	CN_out_sig(154);
VN_in_sig(2084)	<=	CN_out_sig(155);
VN_in_sig(2844)	<=	CN_out_sig(156);
VN_in_sig(3492)	<=	CN_out_sig(157);
VN_in_sig(3996)	<=	CN_out_sig(158);
VN_in_sig(5044)	<=	CN_out_sig(159);
VN_in_sig(124)	<=	CN_out_sig(160);
VN_in_sig(1052)	<=	CN_out_sig(161);
VN_in_sig(1940)	<=	CN_out_sig(162);
VN_in_sig(2088)	<=	CN_out_sig(163);
VN_in_sig(2848)	<=	CN_out_sig(164);
VN_in_sig(3496)	<=	CN_out_sig(165);
VN_in_sig(4000)	<=	CN_out_sig(166);
VN_in_sig(5048)	<=	CN_out_sig(167);
VN_in_sig(128)	<=	CN_out_sig(168);
VN_in_sig(1056)	<=	CN_out_sig(169);
VN_in_sig(1728)	<=	CN_out_sig(170);
VN_in_sig(2092)	<=	CN_out_sig(171);
VN_in_sig(2852)	<=	CN_out_sig(172);
VN_in_sig(3500)	<=	CN_out_sig(173);
VN_in_sig(4004)	<=	CN_out_sig(174);
VN_in_sig(5052)	<=	CN_out_sig(175);
VN_in_sig(132)	<=	CN_out_sig(176);
VN_in_sig(1060)	<=	CN_out_sig(177);
VN_in_sig(1732)	<=	CN_out_sig(178);
VN_in_sig(2096)	<=	CN_out_sig(179);
VN_in_sig(2856)	<=	CN_out_sig(180);
VN_in_sig(3504)	<=	CN_out_sig(181);
VN_in_sig(4008)	<=	CN_out_sig(182);
VN_in_sig(5056)	<=	CN_out_sig(183);
VN_in_sig(136)	<=	CN_out_sig(184);
VN_in_sig(1064)	<=	CN_out_sig(185);
VN_in_sig(1736)	<=	CN_out_sig(186);
VN_in_sig(2100)	<=	CN_out_sig(187);
VN_in_sig(2860)	<=	CN_out_sig(188);
VN_in_sig(3508)	<=	CN_out_sig(189);
VN_in_sig(4012)	<=	CN_out_sig(190);
VN_in_sig(5060)	<=	CN_out_sig(191);
VN_in_sig(140)	<=	CN_out_sig(192);
VN_in_sig(1068)	<=	CN_out_sig(193);
VN_in_sig(1740)	<=	CN_out_sig(194);
VN_in_sig(2104)	<=	CN_out_sig(195);
VN_in_sig(2864)	<=	CN_out_sig(196);
VN_in_sig(3512)	<=	CN_out_sig(197);
VN_in_sig(4016)	<=	CN_out_sig(198);
VN_in_sig(5064)	<=	CN_out_sig(199);
VN_in_sig(144)	<=	CN_out_sig(200);
VN_in_sig(1072)	<=	CN_out_sig(201);
VN_in_sig(1744)	<=	CN_out_sig(202);
VN_in_sig(2108)	<=	CN_out_sig(203);
VN_in_sig(2868)	<=	CN_out_sig(204);
VN_in_sig(3516)	<=	CN_out_sig(205);
VN_in_sig(4020)	<=	CN_out_sig(206);
VN_in_sig(5068)	<=	CN_out_sig(207);
VN_in_sig(148)	<=	CN_out_sig(208);
VN_in_sig(1076)	<=	CN_out_sig(209);
VN_in_sig(1748)	<=	CN_out_sig(210);
VN_in_sig(2112)	<=	CN_out_sig(211);
VN_in_sig(2872)	<=	CN_out_sig(212);
VN_in_sig(3520)	<=	CN_out_sig(213);
VN_in_sig(4024)	<=	CN_out_sig(214);
VN_in_sig(5072)	<=	CN_out_sig(215);
VN_in_sig(152)	<=	CN_out_sig(216);
VN_in_sig(864)	<=	CN_out_sig(217);
VN_in_sig(1752)	<=	CN_out_sig(218);
VN_in_sig(2116)	<=	CN_out_sig(219);
VN_in_sig(2876)	<=	CN_out_sig(220);
VN_in_sig(3524)	<=	CN_out_sig(221);
VN_in_sig(4028)	<=	CN_out_sig(222);
VN_in_sig(5076)	<=	CN_out_sig(223);
VN_in_sig(156)	<=	CN_out_sig(224);
VN_in_sig(868)	<=	CN_out_sig(225);
VN_in_sig(1756)	<=	CN_out_sig(226);
VN_in_sig(2120)	<=	CN_out_sig(227);
VN_in_sig(2880)	<=	CN_out_sig(228);
VN_in_sig(3528)	<=	CN_out_sig(229);
VN_in_sig(4032)	<=	CN_out_sig(230);
VN_in_sig(5080)	<=	CN_out_sig(231);
VN_in_sig(160)	<=	CN_out_sig(232);
VN_in_sig(872)	<=	CN_out_sig(233);
VN_in_sig(1760)	<=	CN_out_sig(234);
VN_in_sig(2124)	<=	CN_out_sig(235);
VN_in_sig(2884)	<=	CN_out_sig(236);
VN_in_sig(3532)	<=	CN_out_sig(237);
VN_in_sig(4036)	<=	CN_out_sig(238);
VN_in_sig(5084)	<=	CN_out_sig(239);
VN_in_sig(164)	<=	CN_out_sig(240);
VN_in_sig(876)	<=	CN_out_sig(241);
VN_in_sig(1764)	<=	CN_out_sig(242);
VN_in_sig(2128)	<=	CN_out_sig(243);
VN_in_sig(2888)	<=	CN_out_sig(244);
VN_in_sig(3536)	<=	CN_out_sig(245);
VN_in_sig(4040)	<=	CN_out_sig(246);
VN_in_sig(5088)	<=	CN_out_sig(247);
VN_in_sig(168)	<=	CN_out_sig(248);
VN_in_sig(880)	<=	CN_out_sig(249);
VN_in_sig(1768)	<=	CN_out_sig(250);
VN_in_sig(2132)	<=	CN_out_sig(251);
VN_in_sig(2892)	<=	CN_out_sig(252);
VN_in_sig(3540)	<=	CN_out_sig(253);
VN_in_sig(4044)	<=	CN_out_sig(254);
VN_in_sig(5092)	<=	CN_out_sig(255);
VN_in_sig(172)	<=	CN_out_sig(256);
VN_in_sig(884)	<=	CN_out_sig(257);
VN_in_sig(1772)	<=	CN_out_sig(258);
VN_in_sig(2136)	<=	CN_out_sig(259);
VN_in_sig(2896)	<=	CN_out_sig(260);
VN_in_sig(3544)	<=	CN_out_sig(261);
VN_in_sig(4048)	<=	CN_out_sig(262);
VN_in_sig(5096)	<=	CN_out_sig(263);
VN_in_sig(176)	<=	CN_out_sig(264);
VN_in_sig(888)	<=	CN_out_sig(265);
VN_in_sig(1776)	<=	CN_out_sig(266);
VN_in_sig(2140)	<=	CN_out_sig(267);
VN_in_sig(2900)	<=	CN_out_sig(268);
VN_in_sig(3548)	<=	CN_out_sig(269);
VN_in_sig(4052)	<=	CN_out_sig(270);
VN_in_sig(5100)	<=	CN_out_sig(271);
VN_in_sig(180)	<=	CN_out_sig(272);
VN_in_sig(892)	<=	CN_out_sig(273);
VN_in_sig(1780)	<=	CN_out_sig(274);
VN_in_sig(2144)	<=	CN_out_sig(275);
VN_in_sig(2904)	<=	CN_out_sig(276);
VN_in_sig(3552)	<=	CN_out_sig(277);
VN_in_sig(4056)	<=	CN_out_sig(278);
VN_in_sig(5104)	<=	CN_out_sig(279);
VN_in_sig(184)	<=	CN_out_sig(280);
VN_in_sig(896)	<=	CN_out_sig(281);
VN_in_sig(1784)	<=	CN_out_sig(282);
VN_in_sig(2148)	<=	CN_out_sig(283);
VN_in_sig(2908)	<=	CN_out_sig(284);
VN_in_sig(3556)	<=	CN_out_sig(285);
VN_in_sig(4060)	<=	CN_out_sig(286);
VN_in_sig(5108)	<=	CN_out_sig(287);
VN_in_sig(188)	<=	CN_out_sig(288);
VN_in_sig(900)	<=	CN_out_sig(289);
VN_in_sig(1788)	<=	CN_out_sig(290);
VN_in_sig(2152)	<=	CN_out_sig(291);
VN_in_sig(2912)	<=	CN_out_sig(292);
VN_in_sig(3560)	<=	CN_out_sig(293);
VN_in_sig(4064)	<=	CN_out_sig(294);
VN_in_sig(5112)	<=	CN_out_sig(295);
VN_in_sig(192)	<=	CN_out_sig(296);
VN_in_sig(904)	<=	CN_out_sig(297);
VN_in_sig(1792)	<=	CN_out_sig(298);
VN_in_sig(2156)	<=	CN_out_sig(299);
VN_in_sig(2916)	<=	CN_out_sig(300);
VN_in_sig(3564)	<=	CN_out_sig(301);
VN_in_sig(4068)	<=	CN_out_sig(302);
VN_in_sig(5116)	<=	CN_out_sig(303);
VN_in_sig(196)	<=	CN_out_sig(304);
VN_in_sig(908)	<=	CN_out_sig(305);
VN_in_sig(1796)	<=	CN_out_sig(306);
VN_in_sig(1944)	<=	CN_out_sig(307);
VN_in_sig(2920)	<=	CN_out_sig(308);
VN_in_sig(3568)	<=	CN_out_sig(309);
VN_in_sig(4072)	<=	CN_out_sig(310);
VN_in_sig(5120)	<=	CN_out_sig(311);
VN_in_sig(200)	<=	CN_out_sig(312);
VN_in_sig(912)	<=	CN_out_sig(313);
VN_in_sig(1800)	<=	CN_out_sig(314);
VN_in_sig(1948)	<=	CN_out_sig(315);
VN_in_sig(2924)	<=	CN_out_sig(316);
VN_in_sig(3572)	<=	CN_out_sig(317);
VN_in_sig(4076)	<=	CN_out_sig(318);
VN_in_sig(5124)	<=	CN_out_sig(319);
VN_in_sig(204)	<=	CN_out_sig(320);
VN_in_sig(916)	<=	CN_out_sig(321);
VN_in_sig(1804)	<=	CN_out_sig(322);
VN_in_sig(1952)	<=	CN_out_sig(323);
VN_in_sig(2928)	<=	CN_out_sig(324);
VN_in_sig(3576)	<=	CN_out_sig(325);
VN_in_sig(4080)	<=	CN_out_sig(326);
VN_in_sig(5128)	<=	CN_out_sig(327);
VN_in_sig(208)	<=	CN_out_sig(328);
VN_in_sig(920)	<=	CN_out_sig(329);
VN_in_sig(1808)	<=	CN_out_sig(330);
VN_in_sig(1956)	<=	CN_out_sig(331);
VN_in_sig(2932)	<=	CN_out_sig(332);
VN_in_sig(3580)	<=	CN_out_sig(333);
VN_in_sig(4084)	<=	CN_out_sig(334);
VN_in_sig(5132)	<=	CN_out_sig(335);
VN_in_sig(212)	<=	CN_out_sig(336);
VN_in_sig(924)	<=	CN_out_sig(337);
VN_in_sig(1812)	<=	CN_out_sig(338);
VN_in_sig(1960)	<=	CN_out_sig(339);
VN_in_sig(2936)	<=	CN_out_sig(340);
VN_in_sig(3584)	<=	CN_out_sig(341);
VN_in_sig(4088)	<=	CN_out_sig(342);
VN_in_sig(5136)	<=	CN_out_sig(343);
VN_in_sig(0)	<=	CN_out_sig(344);
VN_in_sig(928)	<=	CN_out_sig(345);
VN_in_sig(1816)	<=	CN_out_sig(346);
VN_in_sig(1964)	<=	CN_out_sig(347);
VN_in_sig(2940)	<=	CN_out_sig(348);
VN_in_sig(3588)	<=	CN_out_sig(349);
VN_in_sig(4092)	<=	CN_out_sig(350);
VN_in_sig(5140)	<=	CN_out_sig(351);
VN_in_sig(4)	<=	CN_out_sig(352);
VN_in_sig(932)	<=	CN_out_sig(353);
VN_in_sig(1820)	<=	CN_out_sig(354);
VN_in_sig(1968)	<=	CN_out_sig(355);
VN_in_sig(2944)	<=	CN_out_sig(356);
VN_in_sig(3592)	<=	CN_out_sig(357);
VN_in_sig(4096)	<=	CN_out_sig(358);
VN_in_sig(5144)	<=	CN_out_sig(359);
VN_in_sig(8)	<=	CN_out_sig(360);
VN_in_sig(936)	<=	CN_out_sig(361);
VN_in_sig(1824)	<=	CN_out_sig(362);
VN_in_sig(1972)	<=	CN_out_sig(363);
VN_in_sig(2948)	<=	CN_out_sig(364);
VN_in_sig(3596)	<=	CN_out_sig(365);
VN_in_sig(4100)	<=	CN_out_sig(366);
VN_in_sig(5148)	<=	CN_out_sig(367);
VN_in_sig(12)	<=	CN_out_sig(368);
VN_in_sig(940)	<=	CN_out_sig(369);
VN_in_sig(1828)	<=	CN_out_sig(370);
VN_in_sig(1976)	<=	CN_out_sig(371);
VN_in_sig(2952)	<=	CN_out_sig(372);
VN_in_sig(3600)	<=	CN_out_sig(373);
VN_in_sig(3888)	<=	CN_out_sig(374);
VN_in_sig(5152)	<=	CN_out_sig(375);
VN_in_sig(16)	<=	CN_out_sig(376);
VN_in_sig(944)	<=	CN_out_sig(377);
VN_in_sig(1832)	<=	CN_out_sig(378);
VN_in_sig(1980)	<=	CN_out_sig(379);
VN_in_sig(2956)	<=	CN_out_sig(380);
VN_in_sig(3604)	<=	CN_out_sig(381);
VN_in_sig(3892)	<=	CN_out_sig(382);
VN_in_sig(5156)	<=	CN_out_sig(383);
VN_in_sig(20)	<=	CN_out_sig(384);
VN_in_sig(948)	<=	CN_out_sig(385);
VN_in_sig(1836)	<=	CN_out_sig(386);
VN_in_sig(1984)	<=	CN_out_sig(387);
VN_in_sig(2960)	<=	CN_out_sig(388);
VN_in_sig(3608)	<=	CN_out_sig(389);
VN_in_sig(3896)	<=	CN_out_sig(390);
VN_in_sig(5160)	<=	CN_out_sig(391);
VN_in_sig(24)	<=	CN_out_sig(392);
VN_in_sig(952)	<=	CN_out_sig(393);
VN_in_sig(1840)	<=	CN_out_sig(394);
VN_in_sig(1988)	<=	CN_out_sig(395);
VN_in_sig(2964)	<=	CN_out_sig(396);
VN_in_sig(3612)	<=	CN_out_sig(397);
VN_in_sig(3900)	<=	CN_out_sig(398);
VN_in_sig(5164)	<=	CN_out_sig(399);
VN_in_sig(28)	<=	CN_out_sig(400);
VN_in_sig(956)	<=	CN_out_sig(401);
VN_in_sig(1844)	<=	CN_out_sig(402);
VN_in_sig(1992)	<=	CN_out_sig(403);
VN_in_sig(2968)	<=	CN_out_sig(404);
VN_in_sig(3616)	<=	CN_out_sig(405);
VN_in_sig(3904)	<=	CN_out_sig(406);
VN_in_sig(5168)	<=	CN_out_sig(407);
VN_in_sig(32)	<=	CN_out_sig(408);
VN_in_sig(960)	<=	CN_out_sig(409);
VN_in_sig(1848)	<=	CN_out_sig(410);
VN_in_sig(1996)	<=	CN_out_sig(411);
VN_in_sig(2972)	<=	CN_out_sig(412);
VN_in_sig(3620)	<=	CN_out_sig(413);
VN_in_sig(3908)	<=	CN_out_sig(414);
VN_in_sig(5172)	<=	CN_out_sig(415);
VN_in_sig(36)	<=	CN_out_sig(416);
VN_in_sig(964)	<=	CN_out_sig(417);
VN_in_sig(1852)	<=	CN_out_sig(418);
VN_in_sig(2000)	<=	CN_out_sig(419);
VN_in_sig(2976)	<=	CN_out_sig(420);
VN_in_sig(3624)	<=	CN_out_sig(421);
VN_in_sig(3912)	<=	CN_out_sig(422);
VN_in_sig(5176)	<=	CN_out_sig(423);
VN_in_sig(40)	<=	CN_out_sig(424);
VN_in_sig(968)	<=	CN_out_sig(425);
VN_in_sig(1856)	<=	CN_out_sig(426);
VN_in_sig(2004)	<=	CN_out_sig(427);
VN_in_sig(2980)	<=	CN_out_sig(428);
VN_in_sig(3628)	<=	CN_out_sig(429);
VN_in_sig(3916)	<=	CN_out_sig(430);
VN_in_sig(5180)	<=	CN_out_sig(431);
VN_in_sig(316)	<=	CN_out_sig(432);
VN_in_sig(1204)	<=	CN_out_sig(433);
VN_in_sig(1412)	<=	CN_out_sig(434);
VN_in_sig(2276)	<=	CN_out_sig(435);
VN_in_sig(3168)	<=	CN_out_sig(436);
VN_in_sig(3808)	<=	CN_out_sig(437);
VN_in_sig(4164)	<=	CN_out_sig(438);
VN_in_sig(4820)	<=	CN_out_sig(439);
VN_in_sig(320)	<=	CN_out_sig(440);
VN_in_sig(1208)	<=	CN_out_sig(441);
VN_in_sig(1416)	<=	CN_out_sig(442);
VN_in_sig(2280)	<=	CN_out_sig(443);
VN_in_sig(3172)	<=	CN_out_sig(444);
VN_in_sig(3812)	<=	CN_out_sig(445);
VN_in_sig(4168)	<=	CN_out_sig(446);
VN_in_sig(4824)	<=	CN_out_sig(447);
VN_in_sig(324)	<=	CN_out_sig(448);
VN_in_sig(1212)	<=	CN_out_sig(449);
VN_in_sig(1420)	<=	CN_out_sig(450);
VN_in_sig(2284)	<=	CN_out_sig(451);
VN_in_sig(3176)	<=	CN_out_sig(452);
VN_in_sig(3816)	<=	CN_out_sig(453);
VN_in_sig(4172)	<=	CN_out_sig(454);
VN_in_sig(4828)	<=	CN_out_sig(455);
VN_in_sig(328)	<=	CN_out_sig(456);
VN_in_sig(1216)	<=	CN_out_sig(457);
VN_in_sig(1424)	<=	CN_out_sig(458);
VN_in_sig(2288)	<=	CN_out_sig(459);
VN_in_sig(3180)	<=	CN_out_sig(460);
VN_in_sig(3820)	<=	CN_out_sig(461);
VN_in_sig(4176)	<=	CN_out_sig(462);
VN_in_sig(4832)	<=	CN_out_sig(463);
VN_in_sig(332)	<=	CN_out_sig(464);
VN_in_sig(1220)	<=	CN_out_sig(465);
VN_in_sig(1428)	<=	CN_out_sig(466);
VN_in_sig(2292)	<=	CN_out_sig(467);
VN_in_sig(3184)	<=	CN_out_sig(468);
VN_in_sig(3824)	<=	CN_out_sig(469);
VN_in_sig(4180)	<=	CN_out_sig(470);
VN_in_sig(4836)	<=	CN_out_sig(471);
VN_in_sig(336)	<=	CN_out_sig(472);
VN_in_sig(1224)	<=	CN_out_sig(473);
VN_in_sig(1432)	<=	CN_out_sig(474);
VN_in_sig(2296)	<=	CN_out_sig(475);
VN_in_sig(3188)	<=	CN_out_sig(476);
VN_in_sig(3828)	<=	CN_out_sig(477);
VN_in_sig(4184)	<=	CN_out_sig(478);
VN_in_sig(4840)	<=	CN_out_sig(479);
VN_in_sig(340)	<=	CN_out_sig(480);
VN_in_sig(1228)	<=	CN_out_sig(481);
VN_in_sig(1436)	<=	CN_out_sig(482);
VN_in_sig(2300)	<=	CN_out_sig(483);
VN_in_sig(3192)	<=	CN_out_sig(484);
VN_in_sig(3832)	<=	CN_out_sig(485);
VN_in_sig(4188)	<=	CN_out_sig(486);
VN_in_sig(4844)	<=	CN_out_sig(487);
VN_in_sig(344)	<=	CN_out_sig(488);
VN_in_sig(1232)	<=	CN_out_sig(489);
VN_in_sig(1440)	<=	CN_out_sig(490);
VN_in_sig(2304)	<=	CN_out_sig(491);
VN_in_sig(3196)	<=	CN_out_sig(492);
VN_in_sig(3836)	<=	CN_out_sig(493);
VN_in_sig(4192)	<=	CN_out_sig(494);
VN_in_sig(4848)	<=	CN_out_sig(495);
VN_in_sig(348)	<=	CN_out_sig(496);
VN_in_sig(1236)	<=	CN_out_sig(497);
VN_in_sig(1444)	<=	CN_out_sig(498);
VN_in_sig(2308)	<=	CN_out_sig(499);
VN_in_sig(3200)	<=	CN_out_sig(500);
VN_in_sig(3840)	<=	CN_out_sig(501);
VN_in_sig(4196)	<=	CN_out_sig(502);
VN_in_sig(4852)	<=	CN_out_sig(503);
VN_in_sig(352)	<=	CN_out_sig(504);
VN_in_sig(1240)	<=	CN_out_sig(505);
VN_in_sig(1448)	<=	CN_out_sig(506);
VN_in_sig(2312)	<=	CN_out_sig(507);
VN_in_sig(3204)	<=	CN_out_sig(508);
VN_in_sig(3844)	<=	CN_out_sig(509);
VN_in_sig(4200)	<=	CN_out_sig(510);
VN_in_sig(4856)	<=	CN_out_sig(511);
VN_in_sig(356)	<=	CN_out_sig(512);
VN_in_sig(1244)	<=	CN_out_sig(513);
VN_in_sig(1452)	<=	CN_out_sig(514);
VN_in_sig(2316)	<=	CN_out_sig(515);
VN_in_sig(3208)	<=	CN_out_sig(516);
VN_in_sig(3848)	<=	CN_out_sig(517);
VN_in_sig(4204)	<=	CN_out_sig(518);
VN_in_sig(4860)	<=	CN_out_sig(519);
VN_in_sig(360)	<=	CN_out_sig(520);
VN_in_sig(1248)	<=	CN_out_sig(521);
VN_in_sig(1456)	<=	CN_out_sig(522);
VN_in_sig(2320)	<=	CN_out_sig(523);
VN_in_sig(3212)	<=	CN_out_sig(524);
VN_in_sig(3852)	<=	CN_out_sig(525);
VN_in_sig(4208)	<=	CN_out_sig(526);
VN_in_sig(4864)	<=	CN_out_sig(527);
VN_in_sig(364)	<=	CN_out_sig(528);
VN_in_sig(1252)	<=	CN_out_sig(529);
VN_in_sig(1460)	<=	CN_out_sig(530);
VN_in_sig(2324)	<=	CN_out_sig(531);
VN_in_sig(3216)	<=	CN_out_sig(532);
VN_in_sig(3856)	<=	CN_out_sig(533);
VN_in_sig(4212)	<=	CN_out_sig(534);
VN_in_sig(4868)	<=	CN_out_sig(535);
VN_in_sig(368)	<=	CN_out_sig(536);
VN_in_sig(1256)	<=	CN_out_sig(537);
VN_in_sig(1464)	<=	CN_out_sig(538);
VN_in_sig(2328)	<=	CN_out_sig(539);
VN_in_sig(3220)	<=	CN_out_sig(540);
VN_in_sig(3860)	<=	CN_out_sig(541);
VN_in_sig(4216)	<=	CN_out_sig(542);
VN_in_sig(4872)	<=	CN_out_sig(543);
VN_in_sig(372)	<=	CN_out_sig(544);
VN_in_sig(1260)	<=	CN_out_sig(545);
VN_in_sig(1468)	<=	CN_out_sig(546);
VN_in_sig(2332)	<=	CN_out_sig(547);
VN_in_sig(3224)	<=	CN_out_sig(548);
VN_in_sig(3864)	<=	CN_out_sig(549);
VN_in_sig(4220)	<=	CN_out_sig(550);
VN_in_sig(4876)	<=	CN_out_sig(551);
VN_in_sig(376)	<=	CN_out_sig(552);
VN_in_sig(1264)	<=	CN_out_sig(553);
VN_in_sig(1472)	<=	CN_out_sig(554);
VN_in_sig(2336)	<=	CN_out_sig(555);
VN_in_sig(3228)	<=	CN_out_sig(556);
VN_in_sig(3868)	<=	CN_out_sig(557);
VN_in_sig(4224)	<=	CN_out_sig(558);
VN_in_sig(4880)	<=	CN_out_sig(559);
VN_in_sig(380)	<=	CN_out_sig(560);
VN_in_sig(1268)	<=	CN_out_sig(561);
VN_in_sig(1476)	<=	CN_out_sig(562);
VN_in_sig(2340)	<=	CN_out_sig(563);
VN_in_sig(3232)	<=	CN_out_sig(564);
VN_in_sig(3872)	<=	CN_out_sig(565);
VN_in_sig(4228)	<=	CN_out_sig(566);
VN_in_sig(4884)	<=	CN_out_sig(567);
VN_in_sig(384)	<=	CN_out_sig(568);
VN_in_sig(1272)	<=	CN_out_sig(569);
VN_in_sig(1480)	<=	CN_out_sig(570);
VN_in_sig(2344)	<=	CN_out_sig(571);
VN_in_sig(3236)	<=	CN_out_sig(572);
VN_in_sig(3876)	<=	CN_out_sig(573);
VN_in_sig(4232)	<=	CN_out_sig(574);
VN_in_sig(4888)	<=	CN_out_sig(575);
VN_in_sig(388)	<=	CN_out_sig(576);
VN_in_sig(1276)	<=	CN_out_sig(577);
VN_in_sig(1484)	<=	CN_out_sig(578);
VN_in_sig(2348)	<=	CN_out_sig(579);
VN_in_sig(3024)	<=	CN_out_sig(580);
VN_in_sig(3880)	<=	CN_out_sig(581);
VN_in_sig(4236)	<=	CN_out_sig(582);
VN_in_sig(4892)	<=	CN_out_sig(583);
VN_in_sig(392)	<=	CN_out_sig(584);
VN_in_sig(1280)	<=	CN_out_sig(585);
VN_in_sig(1488)	<=	CN_out_sig(586);
VN_in_sig(2352)	<=	CN_out_sig(587);
VN_in_sig(3028)	<=	CN_out_sig(588);
VN_in_sig(3884)	<=	CN_out_sig(589);
VN_in_sig(4240)	<=	CN_out_sig(590);
VN_in_sig(4896)	<=	CN_out_sig(591);
VN_in_sig(396)	<=	CN_out_sig(592);
VN_in_sig(1284)	<=	CN_out_sig(593);
VN_in_sig(1492)	<=	CN_out_sig(594);
VN_in_sig(2356)	<=	CN_out_sig(595);
VN_in_sig(3032)	<=	CN_out_sig(596);
VN_in_sig(3672)	<=	CN_out_sig(597);
VN_in_sig(4244)	<=	CN_out_sig(598);
VN_in_sig(4900)	<=	CN_out_sig(599);
VN_in_sig(400)	<=	CN_out_sig(600);
VN_in_sig(1288)	<=	CN_out_sig(601);
VN_in_sig(1496)	<=	CN_out_sig(602);
VN_in_sig(2360)	<=	CN_out_sig(603);
VN_in_sig(3036)	<=	CN_out_sig(604);
VN_in_sig(3676)	<=	CN_out_sig(605);
VN_in_sig(4248)	<=	CN_out_sig(606);
VN_in_sig(4904)	<=	CN_out_sig(607);
VN_in_sig(404)	<=	CN_out_sig(608);
VN_in_sig(1292)	<=	CN_out_sig(609);
VN_in_sig(1500)	<=	CN_out_sig(610);
VN_in_sig(2364)	<=	CN_out_sig(611);
VN_in_sig(3040)	<=	CN_out_sig(612);
VN_in_sig(3680)	<=	CN_out_sig(613);
VN_in_sig(4252)	<=	CN_out_sig(614);
VN_in_sig(4908)	<=	CN_out_sig(615);
VN_in_sig(408)	<=	CN_out_sig(616);
VN_in_sig(1080)	<=	CN_out_sig(617);
VN_in_sig(1504)	<=	CN_out_sig(618);
VN_in_sig(2368)	<=	CN_out_sig(619);
VN_in_sig(3044)	<=	CN_out_sig(620);
VN_in_sig(3684)	<=	CN_out_sig(621);
VN_in_sig(4256)	<=	CN_out_sig(622);
VN_in_sig(4912)	<=	CN_out_sig(623);
VN_in_sig(412)	<=	CN_out_sig(624);
VN_in_sig(1084)	<=	CN_out_sig(625);
VN_in_sig(1508)	<=	CN_out_sig(626);
VN_in_sig(2372)	<=	CN_out_sig(627);
VN_in_sig(3048)	<=	CN_out_sig(628);
VN_in_sig(3688)	<=	CN_out_sig(629);
VN_in_sig(4260)	<=	CN_out_sig(630);
VN_in_sig(4916)	<=	CN_out_sig(631);
VN_in_sig(416)	<=	CN_out_sig(632);
VN_in_sig(1088)	<=	CN_out_sig(633);
VN_in_sig(1296)	<=	CN_out_sig(634);
VN_in_sig(2160)	<=	CN_out_sig(635);
VN_in_sig(3052)	<=	CN_out_sig(636);
VN_in_sig(3692)	<=	CN_out_sig(637);
VN_in_sig(4264)	<=	CN_out_sig(638);
VN_in_sig(4920)	<=	CN_out_sig(639);
VN_in_sig(420)	<=	CN_out_sig(640);
VN_in_sig(1092)	<=	CN_out_sig(641);
VN_in_sig(1300)	<=	CN_out_sig(642);
VN_in_sig(2164)	<=	CN_out_sig(643);
VN_in_sig(3056)	<=	CN_out_sig(644);
VN_in_sig(3696)	<=	CN_out_sig(645);
VN_in_sig(4268)	<=	CN_out_sig(646);
VN_in_sig(4924)	<=	CN_out_sig(647);
VN_in_sig(424)	<=	CN_out_sig(648);
VN_in_sig(1096)	<=	CN_out_sig(649);
VN_in_sig(1304)	<=	CN_out_sig(650);
VN_in_sig(2168)	<=	CN_out_sig(651);
VN_in_sig(3060)	<=	CN_out_sig(652);
VN_in_sig(3700)	<=	CN_out_sig(653);
VN_in_sig(4272)	<=	CN_out_sig(654);
VN_in_sig(4928)	<=	CN_out_sig(655);
VN_in_sig(428)	<=	CN_out_sig(656);
VN_in_sig(1100)	<=	CN_out_sig(657);
VN_in_sig(1308)	<=	CN_out_sig(658);
VN_in_sig(2172)	<=	CN_out_sig(659);
VN_in_sig(3064)	<=	CN_out_sig(660);
VN_in_sig(3704)	<=	CN_out_sig(661);
VN_in_sig(4276)	<=	CN_out_sig(662);
VN_in_sig(4932)	<=	CN_out_sig(663);
VN_in_sig(216)	<=	CN_out_sig(664);
VN_in_sig(1104)	<=	CN_out_sig(665);
VN_in_sig(1312)	<=	CN_out_sig(666);
VN_in_sig(2176)	<=	CN_out_sig(667);
VN_in_sig(3068)	<=	CN_out_sig(668);
VN_in_sig(3708)	<=	CN_out_sig(669);
VN_in_sig(4280)	<=	CN_out_sig(670);
VN_in_sig(4936)	<=	CN_out_sig(671);
VN_in_sig(220)	<=	CN_out_sig(672);
VN_in_sig(1108)	<=	CN_out_sig(673);
VN_in_sig(1316)	<=	CN_out_sig(674);
VN_in_sig(2180)	<=	CN_out_sig(675);
VN_in_sig(3072)	<=	CN_out_sig(676);
VN_in_sig(3712)	<=	CN_out_sig(677);
VN_in_sig(4284)	<=	CN_out_sig(678);
VN_in_sig(4940)	<=	CN_out_sig(679);
VN_in_sig(224)	<=	CN_out_sig(680);
VN_in_sig(1112)	<=	CN_out_sig(681);
VN_in_sig(1320)	<=	CN_out_sig(682);
VN_in_sig(2184)	<=	CN_out_sig(683);
VN_in_sig(3076)	<=	CN_out_sig(684);
VN_in_sig(3716)	<=	CN_out_sig(685);
VN_in_sig(4288)	<=	CN_out_sig(686);
VN_in_sig(4944)	<=	CN_out_sig(687);
VN_in_sig(228)	<=	CN_out_sig(688);
VN_in_sig(1116)	<=	CN_out_sig(689);
VN_in_sig(1324)	<=	CN_out_sig(690);
VN_in_sig(2188)	<=	CN_out_sig(691);
VN_in_sig(3080)	<=	CN_out_sig(692);
VN_in_sig(3720)	<=	CN_out_sig(693);
VN_in_sig(4292)	<=	CN_out_sig(694);
VN_in_sig(4948)	<=	CN_out_sig(695);
VN_in_sig(232)	<=	CN_out_sig(696);
VN_in_sig(1120)	<=	CN_out_sig(697);
VN_in_sig(1328)	<=	CN_out_sig(698);
VN_in_sig(2192)	<=	CN_out_sig(699);
VN_in_sig(3084)	<=	CN_out_sig(700);
VN_in_sig(3724)	<=	CN_out_sig(701);
VN_in_sig(4296)	<=	CN_out_sig(702);
VN_in_sig(4952)	<=	CN_out_sig(703);
VN_in_sig(236)	<=	CN_out_sig(704);
VN_in_sig(1124)	<=	CN_out_sig(705);
VN_in_sig(1332)	<=	CN_out_sig(706);
VN_in_sig(2196)	<=	CN_out_sig(707);
VN_in_sig(3088)	<=	CN_out_sig(708);
VN_in_sig(3728)	<=	CN_out_sig(709);
VN_in_sig(4300)	<=	CN_out_sig(710);
VN_in_sig(4956)	<=	CN_out_sig(711);
VN_in_sig(240)	<=	CN_out_sig(712);
VN_in_sig(1128)	<=	CN_out_sig(713);
VN_in_sig(1336)	<=	CN_out_sig(714);
VN_in_sig(2200)	<=	CN_out_sig(715);
VN_in_sig(3092)	<=	CN_out_sig(716);
VN_in_sig(3732)	<=	CN_out_sig(717);
VN_in_sig(4304)	<=	CN_out_sig(718);
VN_in_sig(4960)	<=	CN_out_sig(719);
VN_in_sig(244)	<=	CN_out_sig(720);
VN_in_sig(1132)	<=	CN_out_sig(721);
VN_in_sig(1340)	<=	CN_out_sig(722);
VN_in_sig(2204)	<=	CN_out_sig(723);
VN_in_sig(3096)	<=	CN_out_sig(724);
VN_in_sig(3736)	<=	CN_out_sig(725);
VN_in_sig(4308)	<=	CN_out_sig(726);
VN_in_sig(4964)	<=	CN_out_sig(727);
VN_in_sig(248)	<=	CN_out_sig(728);
VN_in_sig(1136)	<=	CN_out_sig(729);
VN_in_sig(1344)	<=	CN_out_sig(730);
VN_in_sig(2208)	<=	CN_out_sig(731);
VN_in_sig(3100)	<=	CN_out_sig(732);
VN_in_sig(3740)	<=	CN_out_sig(733);
VN_in_sig(4312)	<=	CN_out_sig(734);
VN_in_sig(4752)	<=	CN_out_sig(735);
VN_in_sig(252)	<=	CN_out_sig(736);
VN_in_sig(1140)	<=	CN_out_sig(737);
VN_in_sig(1348)	<=	CN_out_sig(738);
VN_in_sig(2212)	<=	CN_out_sig(739);
VN_in_sig(3104)	<=	CN_out_sig(740);
VN_in_sig(3744)	<=	CN_out_sig(741);
VN_in_sig(4316)	<=	CN_out_sig(742);
VN_in_sig(4756)	<=	CN_out_sig(743);
VN_in_sig(256)	<=	CN_out_sig(744);
VN_in_sig(1144)	<=	CN_out_sig(745);
VN_in_sig(1352)	<=	CN_out_sig(746);
VN_in_sig(2216)	<=	CN_out_sig(747);
VN_in_sig(3108)	<=	CN_out_sig(748);
VN_in_sig(3748)	<=	CN_out_sig(749);
VN_in_sig(4104)	<=	CN_out_sig(750);
VN_in_sig(4760)	<=	CN_out_sig(751);
VN_in_sig(260)	<=	CN_out_sig(752);
VN_in_sig(1148)	<=	CN_out_sig(753);
VN_in_sig(1356)	<=	CN_out_sig(754);
VN_in_sig(2220)	<=	CN_out_sig(755);
VN_in_sig(3112)	<=	CN_out_sig(756);
VN_in_sig(3752)	<=	CN_out_sig(757);
VN_in_sig(4108)	<=	CN_out_sig(758);
VN_in_sig(4764)	<=	CN_out_sig(759);
VN_in_sig(264)	<=	CN_out_sig(760);
VN_in_sig(1152)	<=	CN_out_sig(761);
VN_in_sig(1360)	<=	CN_out_sig(762);
VN_in_sig(2224)	<=	CN_out_sig(763);
VN_in_sig(3116)	<=	CN_out_sig(764);
VN_in_sig(3756)	<=	CN_out_sig(765);
VN_in_sig(4112)	<=	CN_out_sig(766);
VN_in_sig(4768)	<=	CN_out_sig(767);
VN_in_sig(268)	<=	CN_out_sig(768);
VN_in_sig(1156)	<=	CN_out_sig(769);
VN_in_sig(1364)	<=	CN_out_sig(770);
VN_in_sig(2228)	<=	CN_out_sig(771);
VN_in_sig(3120)	<=	CN_out_sig(772);
VN_in_sig(3760)	<=	CN_out_sig(773);
VN_in_sig(4116)	<=	CN_out_sig(774);
VN_in_sig(4772)	<=	CN_out_sig(775);
VN_in_sig(272)	<=	CN_out_sig(776);
VN_in_sig(1160)	<=	CN_out_sig(777);
VN_in_sig(1368)	<=	CN_out_sig(778);
VN_in_sig(2232)	<=	CN_out_sig(779);
VN_in_sig(3124)	<=	CN_out_sig(780);
VN_in_sig(3764)	<=	CN_out_sig(781);
VN_in_sig(4120)	<=	CN_out_sig(782);
VN_in_sig(4776)	<=	CN_out_sig(783);
VN_in_sig(276)	<=	CN_out_sig(784);
VN_in_sig(1164)	<=	CN_out_sig(785);
VN_in_sig(1372)	<=	CN_out_sig(786);
VN_in_sig(2236)	<=	CN_out_sig(787);
VN_in_sig(3128)	<=	CN_out_sig(788);
VN_in_sig(3768)	<=	CN_out_sig(789);
VN_in_sig(4124)	<=	CN_out_sig(790);
VN_in_sig(4780)	<=	CN_out_sig(791);
VN_in_sig(280)	<=	CN_out_sig(792);
VN_in_sig(1168)	<=	CN_out_sig(793);
VN_in_sig(1376)	<=	CN_out_sig(794);
VN_in_sig(2240)	<=	CN_out_sig(795);
VN_in_sig(3132)	<=	CN_out_sig(796);
VN_in_sig(3772)	<=	CN_out_sig(797);
VN_in_sig(4128)	<=	CN_out_sig(798);
VN_in_sig(4784)	<=	CN_out_sig(799);
VN_in_sig(284)	<=	CN_out_sig(800);
VN_in_sig(1172)	<=	CN_out_sig(801);
VN_in_sig(1380)	<=	CN_out_sig(802);
VN_in_sig(2244)	<=	CN_out_sig(803);
VN_in_sig(3136)	<=	CN_out_sig(804);
VN_in_sig(3776)	<=	CN_out_sig(805);
VN_in_sig(4132)	<=	CN_out_sig(806);
VN_in_sig(4788)	<=	CN_out_sig(807);
VN_in_sig(288)	<=	CN_out_sig(808);
VN_in_sig(1176)	<=	CN_out_sig(809);
VN_in_sig(1384)	<=	CN_out_sig(810);
VN_in_sig(2248)	<=	CN_out_sig(811);
VN_in_sig(3140)	<=	CN_out_sig(812);
VN_in_sig(3780)	<=	CN_out_sig(813);
VN_in_sig(4136)	<=	CN_out_sig(814);
VN_in_sig(4792)	<=	CN_out_sig(815);
VN_in_sig(292)	<=	CN_out_sig(816);
VN_in_sig(1180)	<=	CN_out_sig(817);
VN_in_sig(1388)	<=	CN_out_sig(818);
VN_in_sig(2252)	<=	CN_out_sig(819);
VN_in_sig(3144)	<=	CN_out_sig(820);
VN_in_sig(3784)	<=	CN_out_sig(821);
VN_in_sig(4140)	<=	CN_out_sig(822);
VN_in_sig(4796)	<=	CN_out_sig(823);
VN_in_sig(296)	<=	CN_out_sig(824);
VN_in_sig(1184)	<=	CN_out_sig(825);
VN_in_sig(1392)	<=	CN_out_sig(826);
VN_in_sig(2256)	<=	CN_out_sig(827);
VN_in_sig(3148)	<=	CN_out_sig(828);
VN_in_sig(3788)	<=	CN_out_sig(829);
VN_in_sig(4144)	<=	CN_out_sig(830);
VN_in_sig(4800)	<=	CN_out_sig(831);
VN_in_sig(300)	<=	CN_out_sig(832);
VN_in_sig(1188)	<=	CN_out_sig(833);
VN_in_sig(1396)	<=	CN_out_sig(834);
VN_in_sig(2260)	<=	CN_out_sig(835);
VN_in_sig(3152)	<=	CN_out_sig(836);
VN_in_sig(3792)	<=	CN_out_sig(837);
VN_in_sig(4148)	<=	CN_out_sig(838);
VN_in_sig(4804)	<=	CN_out_sig(839);
VN_in_sig(304)	<=	CN_out_sig(840);
VN_in_sig(1192)	<=	CN_out_sig(841);
VN_in_sig(1400)	<=	CN_out_sig(842);
VN_in_sig(2264)	<=	CN_out_sig(843);
VN_in_sig(3156)	<=	CN_out_sig(844);
VN_in_sig(3796)	<=	CN_out_sig(845);
VN_in_sig(4152)	<=	CN_out_sig(846);
VN_in_sig(4808)	<=	CN_out_sig(847);
VN_in_sig(308)	<=	CN_out_sig(848);
VN_in_sig(1196)	<=	CN_out_sig(849);
VN_in_sig(1404)	<=	CN_out_sig(850);
VN_in_sig(2268)	<=	CN_out_sig(851);
VN_in_sig(3160)	<=	CN_out_sig(852);
VN_in_sig(3800)	<=	CN_out_sig(853);
VN_in_sig(4156)	<=	CN_out_sig(854);
VN_in_sig(4812)	<=	CN_out_sig(855);
VN_in_sig(312)	<=	CN_out_sig(856);
VN_in_sig(1200)	<=	CN_out_sig(857);
VN_in_sig(1408)	<=	CN_out_sig(858);
VN_in_sig(2272)	<=	CN_out_sig(859);
VN_in_sig(3164)	<=	CN_out_sig(860);
VN_in_sig(3804)	<=	CN_out_sig(861);
VN_in_sig(4160)	<=	CN_out_sig(862);
VN_in_sig(4816)	<=	CN_out_sig(863);
VN_in_sig(608)	<=	CN_out_sig(864);
VN_in_sig(664)	<=	CN_out_sig(865);
VN_in_sig(1556)	<=	CN_out_sig(866);
VN_in_sig(2384)	<=	CN_out_sig(867);
VN_in_sig(2792)	<=	CN_out_sig(868);
VN_in_sig(3448)	<=	CN_out_sig(869);
VN_in_sig(4440)	<=	CN_out_sig(870);
VN_in_sig(4668)	<=	CN_out_sig(871);
VN_in_sig(612)	<=	CN_out_sig(872);
VN_in_sig(668)	<=	CN_out_sig(873);
VN_in_sig(1560)	<=	CN_out_sig(874);
VN_in_sig(2388)	<=	CN_out_sig(875);
VN_in_sig(2796)	<=	CN_out_sig(876);
VN_in_sig(3452)	<=	CN_out_sig(877);
VN_in_sig(4444)	<=	CN_out_sig(878);
VN_in_sig(4672)	<=	CN_out_sig(879);
VN_in_sig(616)	<=	CN_out_sig(880);
VN_in_sig(672)	<=	CN_out_sig(881);
VN_in_sig(1564)	<=	CN_out_sig(882);
VN_in_sig(2392)	<=	CN_out_sig(883);
VN_in_sig(2800)	<=	CN_out_sig(884);
VN_in_sig(3240)	<=	CN_out_sig(885);
VN_in_sig(4448)	<=	CN_out_sig(886);
VN_in_sig(4676)	<=	CN_out_sig(887);
VN_in_sig(620)	<=	CN_out_sig(888);
VN_in_sig(676)	<=	CN_out_sig(889);
VN_in_sig(1568)	<=	CN_out_sig(890);
VN_in_sig(2396)	<=	CN_out_sig(891);
VN_in_sig(2804)	<=	CN_out_sig(892);
VN_in_sig(3244)	<=	CN_out_sig(893);
VN_in_sig(4452)	<=	CN_out_sig(894);
VN_in_sig(4680)	<=	CN_out_sig(895);
VN_in_sig(624)	<=	CN_out_sig(896);
VN_in_sig(680)	<=	CN_out_sig(897);
VN_in_sig(1572)	<=	CN_out_sig(898);
VN_in_sig(2400)	<=	CN_out_sig(899);
VN_in_sig(2592)	<=	CN_out_sig(900);
VN_in_sig(3248)	<=	CN_out_sig(901);
VN_in_sig(4456)	<=	CN_out_sig(902);
VN_in_sig(4684)	<=	CN_out_sig(903);
VN_in_sig(628)	<=	CN_out_sig(904);
VN_in_sig(684)	<=	CN_out_sig(905);
VN_in_sig(1576)	<=	CN_out_sig(906);
VN_in_sig(2404)	<=	CN_out_sig(907);
VN_in_sig(2596)	<=	CN_out_sig(908);
VN_in_sig(3252)	<=	CN_out_sig(909);
VN_in_sig(4460)	<=	CN_out_sig(910);
VN_in_sig(4688)	<=	CN_out_sig(911);
VN_in_sig(632)	<=	CN_out_sig(912);
VN_in_sig(688)	<=	CN_out_sig(913);
VN_in_sig(1580)	<=	CN_out_sig(914);
VN_in_sig(2408)	<=	CN_out_sig(915);
VN_in_sig(2600)	<=	CN_out_sig(916);
VN_in_sig(3256)	<=	CN_out_sig(917);
VN_in_sig(4464)	<=	CN_out_sig(918);
VN_in_sig(4692)	<=	CN_out_sig(919);
VN_in_sig(636)	<=	CN_out_sig(920);
VN_in_sig(692)	<=	CN_out_sig(921);
VN_in_sig(1584)	<=	CN_out_sig(922);
VN_in_sig(2412)	<=	CN_out_sig(923);
VN_in_sig(2604)	<=	CN_out_sig(924);
VN_in_sig(3260)	<=	CN_out_sig(925);
VN_in_sig(4468)	<=	CN_out_sig(926);
VN_in_sig(4696)	<=	CN_out_sig(927);
VN_in_sig(640)	<=	CN_out_sig(928);
VN_in_sig(696)	<=	CN_out_sig(929);
VN_in_sig(1588)	<=	CN_out_sig(930);
VN_in_sig(2416)	<=	CN_out_sig(931);
VN_in_sig(2608)	<=	CN_out_sig(932);
VN_in_sig(3264)	<=	CN_out_sig(933);
VN_in_sig(4472)	<=	CN_out_sig(934);
VN_in_sig(4700)	<=	CN_out_sig(935);
VN_in_sig(644)	<=	CN_out_sig(936);
VN_in_sig(700)	<=	CN_out_sig(937);
VN_in_sig(1592)	<=	CN_out_sig(938);
VN_in_sig(2420)	<=	CN_out_sig(939);
VN_in_sig(2612)	<=	CN_out_sig(940);
VN_in_sig(3268)	<=	CN_out_sig(941);
VN_in_sig(4476)	<=	CN_out_sig(942);
VN_in_sig(4704)	<=	CN_out_sig(943);
VN_in_sig(432)	<=	CN_out_sig(944);
VN_in_sig(704)	<=	CN_out_sig(945);
VN_in_sig(1596)	<=	CN_out_sig(946);
VN_in_sig(2424)	<=	CN_out_sig(947);
VN_in_sig(2616)	<=	CN_out_sig(948);
VN_in_sig(3272)	<=	CN_out_sig(949);
VN_in_sig(4480)	<=	CN_out_sig(950);
VN_in_sig(4708)	<=	CN_out_sig(951);
VN_in_sig(436)	<=	CN_out_sig(952);
VN_in_sig(708)	<=	CN_out_sig(953);
VN_in_sig(1600)	<=	CN_out_sig(954);
VN_in_sig(2428)	<=	CN_out_sig(955);
VN_in_sig(2620)	<=	CN_out_sig(956);
VN_in_sig(3276)	<=	CN_out_sig(957);
VN_in_sig(4484)	<=	CN_out_sig(958);
VN_in_sig(4712)	<=	CN_out_sig(959);
VN_in_sig(440)	<=	CN_out_sig(960);
VN_in_sig(712)	<=	CN_out_sig(961);
VN_in_sig(1604)	<=	CN_out_sig(962);
VN_in_sig(2432)	<=	CN_out_sig(963);
VN_in_sig(2624)	<=	CN_out_sig(964);
VN_in_sig(3280)	<=	CN_out_sig(965);
VN_in_sig(4488)	<=	CN_out_sig(966);
VN_in_sig(4716)	<=	CN_out_sig(967);
VN_in_sig(444)	<=	CN_out_sig(968);
VN_in_sig(716)	<=	CN_out_sig(969);
VN_in_sig(1608)	<=	CN_out_sig(970);
VN_in_sig(2436)	<=	CN_out_sig(971);
VN_in_sig(2628)	<=	CN_out_sig(972);
VN_in_sig(3284)	<=	CN_out_sig(973);
VN_in_sig(4492)	<=	CN_out_sig(974);
VN_in_sig(4720)	<=	CN_out_sig(975);
VN_in_sig(448)	<=	CN_out_sig(976);
VN_in_sig(720)	<=	CN_out_sig(977);
VN_in_sig(1612)	<=	CN_out_sig(978);
VN_in_sig(2440)	<=	CN_out_sig(979);
VN_in_sig(2632)	<=	CN_out_sig(980);
VN_in_sig(3288)	<=	CN_out_sig(981);
VN_in_sig(4496)	<=	CN_out_sig(982);
VN_in_sig(4724)	<=	CN_out_sig(983);
VN_in_sig(452)	<=	CN_out_sig(984);
VN_in_sig(724)	<=	CN_out_sig(985);
VN_in_sig(1616)	<=	CN_out_sig(986);
VN_in_sig(2444)	<=	CN_out_sig(987);
VN_in_sig(2636)	<=	CN_out_sig(988);
VN_in_sig(3292)	<=	CN_out_sig(989);
VN_in_sig(4500)	<=	CN_out_sig(990);
VN_in_sig(4728)	<=	CN_out_sig(991);
VN_in_sig(456)	<=	CN_out_sig(992);
VN_in_sig(728)	<=	CN_out_sig(993);
VN_in_sig(1620)	<=	CN_out_sig(994);
VN_in_sig(2448)	<=	CN_out_sig(995);
VN_in_sig(2640)	<=	CN_out_sig(996);
VN_in_sig(3296)	<=	CN_out_sig(997);
VN_in_sig(4504)	<=	CN_out_sig(998);
VN_in_sig(4732)	<=	CN_out_sig(999);
VN_in_sig(460)	<=	CN_out_sig(1000);
VN_in_sig(732)	<=	CN_out_sig(1001);
VN_in_sig(1624)	<=	CN_out_sig(1002);
VN_in_sig(2452)	<=	CN_out_sig(1003);
VN_in_sig(2644)	<=	CN_out_sig(1004);
VN_in_sig(3300)	<=	CN_out_sig(1005);
VN_in_sig(4508)	<=	CN_out_sig(1006);
VN_in_sig(4736)	<=	CN_out_sig(1007);
VN_in_sig(464)	<=	CN_out_sig(1008);
VN_in_sig(736)	<=	CN_out_sig(1009);
VN_in_sig(1628)	<=	CN_out_sig(1010);
VN_in_sig(2456)	<=	CN_out_sig(1011);
VN_in_sig(2648)	<=	CN_out_sig(1012);
VN_in_sig(3304)	<=	CN_out_sig(1013);
VN_in_sig(4512)	<=	CN_out_sig(1014);
VN_in_sig(4740)	<=	CN_out_sig(1015);
VN_in_sig(468)	<=	CN_out_sig(1016);
VN_in_sig(740)	<=	CN_out_sig(1017);
VN_in_sig(1632)	<=	CN_out_sig(1018);
VN_in_sig(2460)	<=	CN_out_sig(1019);
VN_in_sig(2652)	<=	CN_out_sig(1020);
VN_in_sig(3308)	<=	CN_out_sig(1021);
VN_in_sig(4516)	<=	CN_out_sig(1022);
VN_in_sig(4744)	<=	CN_out_sig(1023);
VN_in_sig(472)	<=	CN_out_sig(1024);
VN_in_sig(744)	<=	CN_out_sig(1025);
VN_in_sig(1636)	<=	CN_out_sig(1026);
VN_in_sig(2464)	<=	CN_out_sig(1027);
VN_in_sig(2656)	<=	CN_out_sig(1028);
VN_in_sig(3312)	<=	CN_out_sig(1029);
VN_in_sig(4520)	<=	CN_out_sig(1030);
VN_in_sig(4748)	<=	CN_out_sig(1031);
VN_in_sig(476)	<=	CN_out_sig(1032);
VN_in_sig(748)	<=	CN_out_sig(1033);
VN_in_sig(1640)	<=	CN_out_sig(1034);
VN_in_sig(2468)	<=	CN_out_sig(1035);
VN_in_sig(2660)	<=	CN_out_sig(1036);
VN_in_sig(3316)	<=	CN_out_sig(1037);
VN_in_sig(4524)	<=	CN_out_sig(1038);
VN_in_sig(4536)	<=	CN_out_sig(1039);
VN_in_sig(480)	<=	CN_out_sig(1040);
VN_in_sig(752)	<=	CN_out_sig(1041);
VN_in_sig(1644)	<=	CN_out_sig(1042);
VN_in_sig(2472)	<=	CN_out_sig(1043);
VN_in_sig(2664)	<=	CN_out_sig(1044);
VN_in_sig(3320)	<=	CN_out_sig(1045);
VN_in_sig(4528)	<=	CN_out_sig(1046);
VN_in_sig(4540)	<=	CN_out_sig(1047);
VN_in_sig(484)	<=	CN_out_sig(1048);
VN_in_sig(756)	<=	CN_out_sig(1049);
VN_in_sig(1648)	<=	CN_out_sig(1050);
VN_in_sig(2476)	<=	CN_out_sig(1051);
VN_in_sig(2668)	<=	CN_out_sig(1052);
VN_in_sig(3324)	<=	CN_out_sig(1053);
VN_in_sig(4532)	<=	CN_out_sig(1054);
VN_in_sig(4544)	<=	CN_out_sig(1055);
VN_in_sig(488)	<=	CN_out_sig(1056);
VN_in_sig(760)	<=	CN_out_sig(1057);
VN_in_sig(1652)	<=	CN_out_sig(1058);
VN_in_sig(2480)	<=	CN_out_sig(1059);
VN_in_sig(2672)	<=	CN_out_sig(1060);
VN_in_sig(3328)	<=	CN_out_sig(1061);
VN_in_sig(4320)	<=	CN_out_sig(1062);
VN_in_sig(4548)	<=	CN_out_sig(1063);
VN_in_sig(492)	<=	CN_out_sig(1064);
VN_in_sig(764)	<=	CN_out_sig(1065);
VN_in_sig(1656)	<=	CN_out_sig(1066);
VN_in_sig(2484)	<=	CN_out_sig(1067);
VN_in_sig(2676)	<=	CN_out_sig(1068);
VN_in_sig(3332)	<=	CN_out_sig(1069);
VN_in_sig(4324)	<=	CN_out_sig(1070);
VN_in_sig(4552)	<=	CN_out_sig(1071);
VN_in_sig(496)	<=	CN_out_sig(1072);
VN_in_sig(768)	<=	CN_out_sig(1073);
VN_in_sig(1660)	<=	CN_out_sig(1074);
VN_in_sig(2488)	<=	CN_out_sig(1075);
VN_in_sig(2680)	<=	CN_out_sig(1076);
VN_in_sig(3336)	<=	CN_out_sig(1077);
VN_in_sig(4328)	<=	CN_out_sig(1078);
VN_in_sig(4556)	<=	CN_out_sig(1079);
VN_in_sig(500)	<=	CN_out_sig(1080);
VN_in_sig(772)	<=	CN_out_sig(1081);
VN_in_sig(1664)	<=	CN_out_sig(1082);
VN_in_sig(2492)	<=	CN_out_sig(1083);
VN_in_sig(2684)	<=	CN_out_sig(1084);
VN_in_sig(3340)	<=	CN_out_sig(1085);
VN_in_sig(4332)	<=	CN_out_sig(1086);
VN_in_sig(4560)	<=	CN_out_sig(1087);
VN_in_sig(504)	<=	CN_out_sig(1088);
VN_in_sig(776)	<=	CN_out_sig(1089);
VN_in_sig(1668)	<=	CN_out_sig(1090);
VN_in_sig(2496)	<=	CN_out_sig(1091);
VN_in_sig(2688)	<=	CN_out_sig(1092);
VN_in_sig(3344)	<=	CN_out_sig(1093);
VN_in_sig(4336)	<=	CN_out_sig(1094);
VN_in_sig(4564)	<=	CN_out_sig(1095);
VN_in_sig(508)	<=	CN_out_sig(1096);
VN_in_sig(780)	<=	CN_out_sig(1097);
VN_in_sig(1672)	<=	CN_out_sig(1098);
VN_in_sig(2500)	<=	CN_out_sig(1099);
VN_in_sig(2692)	<=	CN_out_sig(1100);
VN_in_sig(3348)	<=	CN_out_sig(1101);
VN_in_sig(4340)	<=	CN_out_sig(1102);
VN_in_sig(4568)	<=	CN_out_sig(1103);
VN_in_sig(512)	<=	CN_out_sig(1104);
VN_in_sig(784)	<=	CN_out_sig(1105);
VN_in_sig(1676)	<=	CN_out_sig(1106);
VN_in_sig(2504)	<=	CN_out_sig(1107);
VN_in_sig(2696)	<=	CN_out_sig(1108);
VN_in_sig(3352)	<=	CN_out_sig(1109);
VN_in_sig(4344)	<=	CN_out_sig(1110);
VN_in_sig(4572)	<=	CN_out_sig(1111);
VN_in_sig(516)	<=	CN_out_sig(1112);
VN_in_sig(788)	<=	CN_out_sig(1113);
VN_in_sig(1680)	<=	CN_out_sig(1114);
VN_in_sig(2508)	<=	CN_out_sig(1115);
VN_in_sig(2700)	<=	CN_out_sig(1116);
VN_in_sig(3356)	<=	CN_out_sig(1117);
VN_in_sig(4348)	<=	CN_out_sig(1118);
VN_in_sig(4576)	<=	CN_out_sig(1119);
VN_in_sig(520)	<=	CN_out_sig(1120);
VN_in_sig(792)	<=	CN_out_sig(1121);
VN_in_sig(1684)	<=	CN_out_sig(1122);
VN_in_sig(2512)	<=	CN_out_sig(1123);
VN_in_sig(2704)	<=	CN_out_sig(1124);
VN_in_sig(3360)	<=	CN_out_sig(1125);
VN_in_sig(4352)	<=	CN_out_sig(1126);
VN_in_sig(4580)	<=	CN_out_sig(1127);
VN_in_sig(524)	<=	CN_out_sig(1128);
VN_in_sig(796)	<=	CN_out_sig(1129);
VN_in_sig(1688)	<=	CN_out_sig(1130);
VN_in_sig(2516)	<=	CN_out_sig(1131);
VN_in_sig(2708)	<=	CN_out_sig(1132);
VN_in_sig(3364)	<=	CN_out_sig(1133);
VN_in_sig(4356)	<=	CN_out_sig(1134);
VN_in_sig(4584)	<=	CN_out_sig(1135);
VN_in_sig(528)	<=	CN_out_sig(1136);
VN_in_sig(800)	<=	CN_out_sig(1137);
VN_in_sig(1692)	<=	CN_out_sig(1138);
VN_in_sig(2520)	<=	CN_out_sig(1139);
VN_in_sig(2712)	<=	CN_out_sig(1140);
VN_in_sig(3368)	<=	CN_out_sig(1141);
VN_in_sig(4360)	<=	CN_out_sig(1142);
VN_in_sig(4588)	<=	CN_out_sig(1143);
VN_in_sig(532)	<=	CN_out_sig(1144);
VN_in_sig(804)	<=	CN_out_sig(1145);
VN_in_sig(1696)	<=	CN_out_sig(1146);
VN_in_sig(2524)	<=	CN_out_sig(1147);
VN_in_sig(2716)	<=	CN_out_sig(1148);
VN_in_sig(3372)	<=	CN_out_sig(1149);
VN_in_sig(4364)	<=	CN_out_sig(1150);
VN_in_sig(4592)	<=	CN_out_sig(1151);
VN_in_sig(536)	<=	CN_out_sig(1152);
VN_in_sig(808)	<=	CN_out_sig(1153);
VN_in_sig(1700)	<=	CN_out_sig(1154);
VN_in_sig(2528)	<=	CN_out_sig(1155);
VN_in_sig(2720)	<=	CN_out_sig(1156);
VN_in_sig(3376)	<=	CN_out_sig(1157);
VN_in_sig(4368)	<=	CN_out_sig(1158);
VN_in_sig(4596)	<=	CN_out_sig(1159);
VN_in_sig(540)	<=	CN_out_sig(1160);
VN_in_sig(812)	<=	CN_out_sig(1161);
VN_in_sig(1704)	<=	CN_out_sig(1162);
VN_in_sig(2532)	<=	CN_out_sig(1163);
VN_in_sig(2724)	<=	CN_out_sig(1164);
VN_in_sig(3380)	<=	CN_out_sig(1165);
VN_in_sig(4372)	<=	CN_out_sig(1166);
VN_in_sig(4600)	<=	CN_out_sig(1167);
VN_in_sig(544)	<=	CN_out_sig(1168);
VN_in_sig(816)	<=	CN_out_sig(1169);
VN_in_sig(1708)	<=	CN_out_sig(1170);
VN_in_sig(2536)	<=	CN_out_sig(1171);
VN_in_sig(2728)	<=	CN_out_sig(1172);
VN_in_sig(3384)	<=	CN_out_sig(1173);
VN_in_sig(4376)	<=	CN_out_sig(1174);
VN_in_sig(4604)	<=	CN_out_sig(1175);
VN_in_sig(548)	<=	CN_out_sig(1176);
VN_in_sig(820)	<=	CN_out_sig(1177);
VN_in_sig(1712)	<=	CN_out_sig(1178);
VN_in_sig(2540)	<=	CN_out_sig(1179);
VN_in_sig(2732)	<=	CN_out_sig(1180);
VN_in_sig(3388)	<=	CN_out_sig(1181);
VN_in_sig(4380)	<=	CN_out_sig(1182);
VN_in_sig(4608)	<=	CN_out_sig(1183);
VN_in_sig(552)	<=	CN_out_sig(1184);
VN_in_sig(824)	<=	CN_out_sig(1185);
VN_in_sig(1716)	<=	CN_out_sig(1186);
VN_in_sig(2544)	<=	CN_out_sig(1187);
VN_in_sig(2736)	<=	CN_out_sig(1188);
VN_in_sig(3392)	<=	CN_out_sig(1189);
VN_in_sig(4384)	<=	CN_out_sig(1190);
VN_in_sig(4612)	<=	CN_out_sig(1191);
VN_in_sig(556)	<=	CN_out_sig(1192);
VN_in_sig(828)	<=	CN_out_sig(1193);
VN_in_sig(1720)	<=	CN_out_sig(1194);
VN_in_sig(2548)	<=	CN_out_sig(1195);
VN_in_sig(2740)	<=	CN_out_sig(1196);
VN_in_sig(3396)	<=	CN_out_sig(1197);
VN_in_sig(4388)	<=	CN_out_sig(1198);
VN_in_sig(4616)	<=	CN_out_sig(1199);
VN_in_sig(560)	<=	CN_out_sig(1200);
VN_in_sig(832)	<=	CN_out_sig(1201);
VN_in_sig(1724)	<=	CN_out_sig(1202);
VN_in_sig(2552)	<=	CN_out_sig(1203);
VN_in_sig(2744)	<=	CN_out_sig(1204);
VN_in_sig(3400)	<=	CN_out_sig(1205);
VN_in_sig(4392)	<=	CN_out_sig(1206);
VN_in_sig(4620)	<=	CN_out_sig(1207);
VN_in_sig(564)	<=	CN_out_sig(1208);
VN_in_sig(836)	<=	CN_out_sig(1209);
VN_in_sig(1512)	<=	CN_out_sig(1210);
VN_in_sig(2556)	<=	CN_out_sig(1211);
VN_in_sig(2748)	<=	CN_out_sig(1212);
VN_in_sig(3404)	<=	CN_out_sig(1213);
VN_in_sig(4396)	<=	CN_out_sig(1214);
VN_in_sig(4624)	<=	CN_out_sig(1215);
VN_in_sig(568)	<=	CN_out_sig(1216);
VN_in_sig(840)	<=	CN_out_sig(1217);
VN_in_sig(1516)	<=	CN_out_sig(1218);
VN_in_sig(2560)	<=	CN_out_sig(1219);
VN_in_sig(2752)	<=	CN_out_sig(1220);
VN_in_sig(3408)	<=	CN_out_sig(1221);
VN_in_sig(4400)	<=	CN_out_sig(1222);
VN_in_sig(4628)	<=	CN_out_sig(1223);
VN_in_sig(572)	<=	CN_out_sig(1224);
VN_in_sig(844)	<=	CN_out_sig(1225);
VN_in_sig(1520)	<=	CN_out_sig(1226);
VN_in_sig(2564)	<=	CN_out_sig(1227);
VN_in_sig(2756)	<=	CN_out_sig(1228);
VN_in_sig(3412)	<=	CN_out_sig(1229);
VN_in_sig(4404)	<=	CN_out_sig(1230);
VN_in_sig(4632)	<=	CN_out_sig(1231);
VN_in_sig(576)	<=	CN_out_sig(1232);
VN_in_sig(848)	<=	CN_out_sig(1233);
VN_in_sig(1524)	<=	CN_out_sig(1234);
VN_in_sig(2568)	<=	CN_out_sig(1235);
VN_in_sig(2760)	<=	CN_out_sig(1236);
VN_in_sig(3416)	<=	CN_out_sig(1237);
VN_in_sig(4408)	<=	CN_out_sig(1238);
VN_in_sig(4636)	<=	CN_out_sig(1239);
VN_in_sig(580)	<=	CN_out_sig(1240);
VN_in_sig(852)	<=	CN_out_sig(1241);
VN_in_sig(1528)	<=	CN_out_sig(1242);
VN_in_sig(2572)	<=	CN_out_sig(1243);
VN_in_sig(2764)	<=	CN_out_sig(1244);
VN_in_sig(3420)	<=	CN_out_sig(1245);
VN_in_sig(4412)	<=	CN_out_sig(1246);
VN_in_sig(4640)	<=	CN_out_sig(1247);
VN_in_sig(584)	<=	CN_out_sig(1248);
VN_in_sig(856)	<=	CN_out_sig(1249);
VN_in_sig(1532)	<=	CN_out_sig(1250);
VN_in_sig(2576)	<=	CN_out_sig(1251);
VN_in_sig(2768)	<=	CN_out_sig(1252);
VN_in_sig(3424)	<=	CN_out_sig(1253);
VN_in_sig(4416)	<=	CN_out_sig(1254);
VN_in_sig(4644)	<=	CN_out_sig(1255);
VN_in_sig(588)	<=	CN_out_sig(1256);
VN_in_sig(860)	<=	CN_out_sig(1257);
VN_in_sig(1536)	<=	CN_out_sig(1258);
VN_in_sig(2580)	<=	CN_out_sig(1259);
VN_in_sig(2772)	<=	CN_out_sig(1260);
VN_in_sig(3428)	<=	CN_out_sig(1261);
VN_in_sig(4420)	<=	CN_out_sig(1262);
VN_in_sig(4648)	<=	CN_out_sig(1263);
VN_in_sig(592)	<=	CN_out_sig(1264);
VN_in_sig(648)	<=	CN_out_sig(1265);
VN_in_sig(1540)	<=	CN_out_sig(1266);
VN_in_sig(2584)	<=	CN_out_sig(1267);
VN_in_sig(2776)	<=	CN_out_sig(1268);
VN_in_sig(3432)	<=	CN_out_sig(1269);
VN_in_sig(4424)	<=	CN_out_sig(1270);
VN_in_sig(4652)	<=	CN_out_sig(1271);
VN_in_sig(596)	<=	CN_out_sig(1272);
VN_in_sig(652)	<=	CN_out_sig(1273);
VN_in_sig(1544)	<=	CN_out_sig(1274);
VN_in_sig(2588)	<=	CN_out_sig(1275);
VN_in_sig(2780)	<=	CN_out_sig(1276);
VN_in_sig(3436)	<=	CN_out_sig(1277);
VN_in_sig(4428)	<=	CN_out_sig(1278);
VN_in_sig(4656)	<=	CN_out_sig(1279);
VN_in_sig(600)	<=	CN_out_sig(1280);
VN_in_sig(656)	<=	CN_out_sig(1281);
VN_in_sig(1548)	<=	CN_out_sig(1282);
VN_in_sig(2376)	<=	CN_out_sig(1283);
VN_in_sig(2784)	<=	CN_out_sig(1284);
VN_in_sig(3440)	<=	CN_out_sig(1285);
VN_in_sig(4432)	<=	CN_out_sig(1286);
VN_in_sig(4660)	<=	CN_out_sig(1287);
VN_in_sig(604)	<=	CN_out_sig(1288);
VN_in_sig(660)	<=	CN_out_sig(1289);
VN_in_sig(1552)	<=	CN_out_sig(1290);
VN_in_sig(2380)	<=	CN_out_sig(1291);
VN_in_sig(2788)	<=	CN_out_sig(1292);
VN_in_sig(3444)	<=	CN_out_sig(1293);
VN_in_sig(4436)	<=	CN_out_sig(1294);
VN_in_sig(4664)	<=	CN_out_sig(1295);
VN_in_sig(109)	<=	CN_out_sig(1296);
VN_in_sig(1001)	<=	CN_out_sig(1297);
VN_in_sig(1377)	<=	CN_out_sig(1298);
VN_in_sig(2025)	<=	CN_out_sig(1299);
VN_in_sig(2861)	<=	CN_out_sig(1300);
VN_in_sig(3565)	<=	CN_out_sig(1301);
VN_in_sig(3905)	<=	CN_out_sig(1302);
VN_in_sig(5077)	<=	CN_out_sig(1303);
VN_in_sig(113)	<=	CN_out_sig(1304);
VN_in_sig(1005)	<=	CN_out_sig(1305);
VN_in_sig(1381)	<=	CN_out_sig(1306);
VN_in_sig(2029)	<=	CN_out_sig(1307);
VN_in_sig(2865)	<=	CN_out_sig(1308);
VN_in_sig(3569)	<=	CN_out_sig(1309);
VN_in_sig(3909)	<=	CN_out_sig(1310);
VN_in_sig(5081)	<=	CN_out_sig(1311);
VN_in_sig(117)	<=	CN_out_sig(1312);
VN_in_sig(1009)	<=	CN_out_sig(1313);
VN_in_sig(1385)	<=	CN_out_sig(1314);
VN_in_sig(2033)	<=	CN_out_sig(1315);
VN_in_sig(2869)	<=	CN_out_sig(1316);
VN_in_sig(3573)	<=	CN_out_sig(1317);
VN_in_sig(3913)	<=	CN_out_sig(1318);
VN_in_sig(5085)	<=	CN_out_sig(1319);
VN_in_sig(121)	<=	CN_out_sig(1320);
VN_in_sig(1013)	<=	CN_out_sig(1321);
VN_in_sig(1389)	<=	CN_out_sig(1322);
VN_in_sig(2037)	<=	CN_out_sig(1323);
VN_in_sig(2873)	<=	CN_out_sig(1324);
VN_in_sig(3577)	<=	CN_out_sig(1325);
VN_in_sig(3917)	<=	CN_out_sig(1326);
VN_in_sig(5089)	<=	CN_out_sig(1327);
VN_in_sig(125)	<=	CN_out_sig(1328);
VN_in_sig(1017)	<=	CN_out_sig(1329);
VN_in_sig(1393)	<=	CN_out_sig(1330);
VN_in_sig(2041)	<=	CN_out_sig(1331);
VN_in_sig(2877)	<=	CN_out_sig(1332);
VN_in_sig(3581)	<=	CN_out_sig(1333);
VN_in_sig(3921)	<=	CN_out_sig(1334);
VN_in_sig(5093)	<=	CN_out_sig(1335);
VN_in_sig(129)	<=	CN_out_sig(1336);
VN_in_sig(1021)	<=	CN_out_sig(1337);
VN_in_sig(1397)	<=	CN_out_sig(1338);
VN_in_sig(2045)	<=	CN_out_sig(1339);
VN_in_sig(2881)	<=	CN_out_sig(1340);
VN_in_sig(3585)	<=	CN_out_sig(1341);
VN_in_sig(3925)	<=	CN_out_sig(1342);
VN_in_sig(5097)	<=	CN_out_sig(1343);
VN_in_sig(133)	<=	CN_out_sig(1344);
VN_in_sig(1025)	<=	CN_out_sig(1345);
VN_in_sig(1401)	<=	CN_out_sig(1346);
VN_in_sig(2049)	<=	CN_out_sig(1347);
VN_in_sig(2885)	<=	CN_out_sig(1348);
VN_in_sig(3589)	<=	CN_out_sig(1349);
VN_in_sig(3929)	<=	CN_out_sig(1350);
VN_in_sig(5101)	<=	CN_out_sig(1351);
VN_in_sig(137)	<=	CN_out_sig(1352);
VN_in_sig(1029)	<=	CN_out_sig(1353);
VN_in_sig(1405)	<=	CN_out_sig(1354);
VN_in_sig(2053)	<=	CN_out_sig(1355);
VN_in_sig(2889)	<=	CN_out_sig(1356);
VN_in_sig(3593)	<=	CN_out_sig(1357);
VN_in_sig(3933)	<=	CN_out_sig(1358);
VN_in_sig(5105)	<=	CN_out_sig(1359);
VN_in_sig(141)	<=	CN_out_sig(1360);
VN_in_sig(1033)	<=	CN_out_sig(1361);
VN_in_sig(1409)	<=	CN_out_sig(1362);
VN_in_sig(2057)	<=	CN_out_sig(1363);
VN_in_sig(2893)	<=	CN_out_sig(1364);
VN_in_sig(3597)	<=	CN_out_sig(1365);
VN_in_sig(3937)	<=	CN_out_sig(1366);
VN_in_sig(5109)	<=	CN_out_sig(1367);
VN_in_sig(145)	<=	CN_out_sig(1368);
VN_in_sig(1037)	<=	CN_out_sig(1369);
VN_in_sig(1413)	<=	CN_out_sig(1370);
VN_in_sig(2061)	<=	CN_out_sig(1371);
VN_in_sig(2897)	<=	CN_out_sig(1372);
VN_in_sig(3601)	<=	CN_out_sig(1373);
VN_in_sig(3941)	<=	CN_out_sig(1374);
VN_in_sig(5113)	<=	CN_out_sig(1375);
VN_in_sig(149)	<=	CN_out_sig(1376);
VN_in_sig(1041)	<=	CN_out_sig(1377);
VN_in_sig(1417)	<=	CN_out_sig(1378);
VN_in_sig(2065)	<=	CN_out_sig(1379);
VN_in_sig(2901)	<=	CN_out_sig(1380);
VN_in_sig(3605)	<=	CN_out_sig(1381);
VN_in_sig(3945)	<=	CN_out_sig(1382);
VN_in_sig(5117)	<=	CN_out_sig(1383);
VN_in_sig(153)	<=	CN_out_sig(1384);
VN_in_sig(1045)	<=	CN_out_sig(1385);
VN_in_sig(1421)	<=	CN_out_sig(1386);
VN_in_sig(2069)	<=	CN_out_sig(1387);
VN_in_sig(2905)	<=	CN_out_sig(1388);
VN_in_sig(3609)	<=	CN_out_sig(1389);
VN_in_sig(3949)	<=	CN_out_sig(1390);
VN_in_sig(5121)	<=	CN_out_sig(1391);
VN_in_sig(157)	<=	CN_out_sig(1392);
VN_in_sig(1049)	<=	CN_out_sig(1393);
VN_in_sig(1425)	<=	CN_out_sig(1394);
VN_in_sig(2073)	<=	CN_out_sig(1395);
VN_in_sig(2909)	<=	CN_out_sig(1396);
VN_in_sig(3613)	<=	CN_out_sig(1397);
VN_in_sig(3953)	<=	CN_out_sig(1398);
VN_in_sig(5125)	<=	CN_out_sig(1399);
VN_in_sig(161)	<=	CN_out_sig(1400);
VN_in_sig(1053)	<=	CN_out_sig(1401);
VN_in_sig(1429)	<=	CN_out_sig(1402);
VN_in_sig(2077)	<=	CN_out_sig(1403);
VN_in_sig(2913)	<=	CN_out_sig(1404);
VN_in_sig(3617)	<=	CN_out_sig(1405);
VN_in_sig(3957)	<=	CN_out_sig(1406);
VN_in_sig(5129)	<=	CN_out_sig(1407);
VN_in_sig(165)	<=	CN_out_sig(1408);
VN_in_sig(1057)	<=	CN_out_sig(1409);
VN_in_sig(1433)	<=	CN_out_sig(1410);
VN_in_sig(2081)	<=	CN_out_sig(1411);
VN_in_sig(2917)	<=	CN_out_sig(1412);
VN_in_sig(3621)	<=	CN_out_sig(1413);
VN_in_sig(3961)	<=	CN_out_sig(1414);
VN_in_sig(5133)	<=	CN_out_sig(1415);
VN_in_sig(169)	<=	CN_out_sig(1416);
VN_in_sig(1061)	<=	CN_out_sig(1417);
VN_in_sig(1437)	<=	CN_out_sig(1418);
VN_in_sig(2085)	<=	CN_out_sig(1419);
VN_in_sig(2921)	<=	CN_out_sig(1420);
VN_in_sig(3625)	<=	CN_out_sig(1421);
VN_in_sig(3965)	<=	CN_out_sig(1422);
VN_in_sig(5137)	<=	CN_out_sig(1423);
VN_in_sig(173)	<=	CN_out_sig(1424);
VN_in_sig(1065)	<=	CN_out_sig(1425);
VN_in_sig(1441)	<=	CN_out_sig(1426);
VN_in_sig(2089)	<=	CN_out_sig(1427);
VN_in_sig(2925)	<=	CN_out_sig(1428);
VN_in_sig(3629)	<=	CN_out_sig(1429);
VN_in_sig(3969)	<=	CN_out_sig(1430);
VN_in_sig(5141)	<=	CN_out_sig(1431);
VN_in_sig(177)	<=	CN_out_sig(1432);
VN_in_sig(1069)	<=	CN_out_sig(1433);
VN_in_sig(1445)	<=	CN_out_sig(1434);
VN_in_sig(2093)	<=	CN_out_sig(1435);
VN_in_sig(2929)	<=	CN_out_sig(1436);
VN_in_sig(3633)	<=	CN_out_sig(1437);
VN_in_sig(3973)	<=	CN_out_sig(1438);
VN_in_sig(5145)	<=	CN_out_sig(1439);
VN_in_sig(181)	<=	CN_out_sig(1440);
VN_in_sig(1073)	<=	CN_out_sig(1441);
VN_in_sig(1449)	<=	CN_out_sig(1442);
VN_in_sig(2097)	<=	CN_out_sig(1443);
VN_in_sig(2933)	<=	CN_out_sig(1444);
VN_in_sig(3637)	<=	CN_out_sig(1445);
VN_in_sig(3977)	<=	CN_out_sig(1446);
VN_in_sig(5149)	<=	CN_out_sig(1447);
VN_in_sig(185)	<=	CN_out_sig(1448);
VN_in_sig(1077)	<=	CN_out_sig(1449);
VN_in_sig(1453)	<=	CN_out_sig(1450);
VN_in_sig(2101)	<=	CN_out_sig(1451);
VN_in_sig(2937)	<=	CN_out_sig(1452);
VN_in_sig(3641)	<=	CN_out_sig(1453);
VN_in_sig(3981)	<=	CN_out_sig(1454);
VN_in_sig(5153)	<=	CN_out_sig(1455);
VN_in_sig(189)	<=	CN_out_sig(1456);
VN_in_sig(865)	<=	CN_out_sig(1457);
VN_in_sig(1457)	<=	CN_out_sig(1458);
VN_in_sig(2105)	<=	CN_out_sig(1459);
VN_in_sig(2941)	<=	CN_out_sig(1460);
VN_in_sig(3645)	<=	CN_out_sig(1461);
VN_in_sig(3985)	<=	CN_out_sig(1462);
VN_in_sig(5157)	<=	CN_out_sig(1463);
VN_in_sig(193)	<=	CN_out_sig(1464);
VN_in_sig(869)	<=	CN_out_sig(1465);
VN_in_sig(1461)	<=	CN_out_sig(1466);
VN_in_sig(2109)	<=	CN_out_sig(1467);
VN_in_sig(2945)	<=	CN_out_sig(1468);
VN_in_sig(3649)	<=	CN_out_sig(1469);
VN_in_sig(3989)	<=	CN_out_sig(1470);
VN_in_sig(5161)	<=	CN_out_sig(1471);
VN_in_sig(197)	<=	CN_out_sig(1472);
VN_in_sig(873)	<=	CN_out_sig(1473);
VN_in_sig(1465)	<=	CN_out_sig(1474);
VN_in_sig(2113)	<=	CN_out_sig(1475);
VN_in_sig(2949)	<=	CN_out_sig(1476);
VN_in_sig(3653)	<=	CN_out_sig(1477);
VN_in_sig(3993)	<=	CN_out_sig(1478);
VN_in_sig(5165)	<=	CN_out_sig(1479);
VN_in_sig(201)	<=	CN_out_sig(1480);
VN_in_sig(877)	<=	CN_out_sig(1481);
VN_in_sig(1469)	<=	CN_out_sig(1482);
VN_in_sig(2117)	<=	CN_out_sig(1483);
VN_in_sig(2953)	<=	CN_out_sig(1484);
VN_in_sig(3657)	<=	CN_out_sig(1485);
VN_in_sig(3997)	<=	CN_out_sig(1486);
VN_in_sig(5169)	<=	CN_out_sig(1487);
VN_in_sig(205)	<=	CN_out_sig(1488);
VN_in_sig(881)	<=	CN_out_sig(1489);
VN_in_sig(1473)	<=	CN_out_sig(1490);
VN_in_sig(2121)	<=	CN_out_sig(1491);
VN_in_sig(2957)	<=	CN_out_sig(1492);
VN_in_sig(3661)	<=	CN_out_sig(1493);
VN_in_sig(4001)	<=	CN_out_sig(1494);
VN_in_sig(5173)	<=	CN_out_sig(1495);
VN_in_sig(209)	<=	CN_out_sig(1496);
VN_in_sig(885)	<=	CN_out_sig(1497);
VN_in_sig(1477)	<=	CN_out_sig(1498);
VN_in_sig(2125)	<=	CN_out_sig(1499);
VN_in_sig(2961)	<=	CN_out_sig(1500);
VN_in_sig(3665)	<=	CN_out_sig(1501);
VN_in_sig(4005)	<=	CN_out_sig(1502);
VN_in_sig(5177)	<=	CN_out_sig(1503);
VN_in_sig(213)	<=	CN_out_sig(1504);
VN_in_sig(889)	<=	CN_out_sig(1505);
VN_in_sig(1481)	<=	CN_out_sig(1506);
VN_in_sig(2129)	<=	CN_out_sig(1507);
VN_in_sig(2965)	<=	CN_out_sig(1508);
VN_in_sig(3669)	<=	CN_out_sig(1509);
VN_in_sig(4009)	<=	CN_out_sig(1510);
VN_in_sig(5181)	<=	CN_out_sig(1511);
VN_in_sig(1)	<=	CN_out_sig(1512);
VN_in_sig(893)	<=	CN_out_sig(1513);
VN_in_sig(1485)	<=	CN_out_sig(1514);
VN_in_sig(2133)	<=	CN_out_sig(1515);
VN_in_sig(2969)	<=	CN_out_sig(1516);
VN_in_sig(3457)	<=	CN_out_sig(1517);
VN_in_sig(4013)	<=	CN_out_sig(1518);
VN_in_sig(4969)	<=	CN_out_sig(1519);
VN_in_sig(5)	<=	CN_out_sig(1520);
VN_in_sig(897)	<=	CN_out_sig(1521);
VN_in_sig(1489)	<=	CN_out_sig(1522);
VN_in_sig(2137)	<=	CN_out_sig(1523);
VN_in_sig(2973)	<=	CN_out_sig(1524);
VN_in_sig(3461)	<=	CN_out_sig(1525);
VN_in_sig(4017)	<=	CN_out_sig(1526);
VN_in_sig(4973)	<=	CN_out_sig(1527);
VN_in_sig(9)	<=	CN_out_sig(1528);
VN_in_sig(901)	<=	CN_out_sig(1529);
VN_in_sig(1493)	<=	CN_out_sig(1530);
VN_in_sig(2141)	<=	CN_out_sig(1531);
VN_in_sig(2977)	<=	CN_out_sig(1532);
VN_in_sig(3465)	<=	CN_out_sig(1533);
VN_in_sig(4021)	<=	CN_out_sig(1534);
VN_in_sig(4977)	<=	CN_out_sig(1535);
VN_in_sig(13)	<=	CN_out_sig(1536);
VN_in_sig(905)	<=	CN_out_sig(1537);
VN_in_sig(1497)	<=	CN_out_sig(1538);
VN_in_sig(2145)	<=	CN_out_sig(1539);
VN_in_sig(2981)	<=	CN_out_sig(1540);
VN_in_sig(3469)	<=	CN_out_sig(1541);
VN_in_sig(4025)	<=	CN_out_sig(1542);
VN_in_sig(4981)	<=	CN_out_sig(1543);
VN_in_sig(17)	<=	CN_out_sig(1544);
VN_in_sig(909)	<=	CN_out_sig(1545);
VN_in_sig(1501)	<=	CN_out_sig(1546);
VN_in_sig(2149)	<=	CN_out_sig(1547);
VN_in_sig(2985)	<=	CN_out_sig(1548);
VN_in_sig(3473)	<=	CN_out_sig(1549);
VN_in_sig(4029)	<=	CN_out_sig(1550);
VN_in_sig(4985)	<=	CN_out_sig(1551);
VN_in_sig(21)	<=	CN_out_sig(1552);
VN_in_sig(913)	<=	CN_out_sig(1553);
VN_in_sig(1505)	<=	CN_out_sig(1554);
VN_in_sig(2153)	<=	CN_out_sig(1555);
VN_in_sig(2989)	<=	CN_out_sig(1556);
VN_in_sig(3477)	<=	CN_out_sig(1557);
VN_in_sig(4033)	<=	CN_out_sig(1558);
VN_in_sig(4989)	<=	CN_out_sig(1559);
VN_in_sig(25)	<=	CN_out_sig(1560);
VN_in_sig(917)	<=	CN_out_sig(1561);
VN_in_sig(1509)	<=	CN_out_sig(1562);
VN_in_sig(2157)	<=	CN_out_sig(1563);
VN_in_sig(2993)	<=	CN_out_sig(1564);
VN_in_sig(3481)	<=	CN_out_sig(1565);
VN_in_sig(4037)	<=	CN_out_sig(1566);
VN_in_sig(4993)	<=	CN_out_sig(1567);
VN_in_sig(29)	<=	CN_out_sig(1568);
VN_in_sig(921)	<=	CN_out_sig(1569);
VN_in_sig(1297)	<=	CN_out_sig(1570);
VN_in_sig(1945)	<=	CN_out_sig(1571);
VN_in_sig(2997)	<=	CN_out_sig(1572);
VN_in_sig(3485)	<=	CN_out_sig(1573);
VN_in_sig(4041)	<=	CN_out_sig(1574);
VN_in_sig(4997)	<=	CN_out_sig(1575);
VN_in_sig(33)	<=	CN_out_sig(1576);
VN_in_sig(925)	<=	CN_out_sig(1577);
VN_in_sig(1301)	<=	CN_out_sig(1578);
VN_in_sig(1949)	<=	CN_out_sig(1579);
VN_in_sig(3001)	<=	CN_out_sig(1580);
VN_in_sig(3489)	<=	CN_out_sig(1581);
VN_in_sig(4045)	<=	CN_out_sig(1582);
VN_in_sig(5001)	<=	CN_out_sig(1583);
VN_in_sig(37)	<=	CN_out_sig(1584);
VN_in_sig(929)	<=	CN_out_sig(1585);
VN_in_sig(1305)	<=	CN_out_sig(1586);
VN_in_sig(1953)	<=	CN_out_sig(1587);
VN_in_sig(3005)	<=	CN_out_sig(1588);
VN_in_sig(3493)	<=	CN_out_sig(1589);
VN_in_sig(4049)	<=	CN_out_sig(1590);
VN_in_sig(5005)	<=	CN_out_sig(1591);
VN_in_sig(41)	<=	CN_out_sig(1592);
VN_in_sig(933)	<=	CN_out_sig(1593);
VN_in_sig(1309)	<=	CN_out_sig(1594);
VN_in_sig(1957)	<=	CN_out_sig(1595);
VN_in_sig(3009)	<=	CN_out_sig(1596);
VN_in_sig(3497)	<=	CN_out_sig(1597);
VN_in_sig(4053)	<=	CN_out_sig(1598);
VN_in_sig(5009)	<=	CN_out_sig(1599);
VN_in_sig(45)	<=	CN_out_sig(1600);
VN_in_sig(937)	<=	CN_out_sig(1601);
VN_in_sig(1313)	<=	CN_out_sig(1602);
VN_in_sig(1961)	<=	CN_out_sig(1603);
VN_in_sig(3013)	<=	CN_out_sig(1604);
VN_in_sig(3501)	<=	CN_out_sig(1605);
VN_in_sig(4057)	<=	CN_out_sig(1606);
VN_in_sig(5013)	<=	CN_out_sig(1607);
VN_in_sig(49)	<=	CN_out_sig(1608);
VN_in_sig(941)	<=	CN_out_sig(1609);
VN_in_sig(1317)	<=	CN_out_sig(1610);
VN_in_sig(1965)	<=	CN_out_sig(1611);
VN_in_sig(3017)	<=	CN_out_sig(1612);
VN_in_sig(3505)	<=	CN_out_sig(1613);
VN_in_sig(4061)	<=	CN_out_sig(1614);
VN_in_sig(5017)	<=	CN_out_sig(1615);
VN_in_sig(53)	<=	CN_out_sig(1616);
VN_in_sig(945)	<=	CN_out_sig(1617);
VN_in_sig(1321)	<=	CN_out_sig(1618);
VN_in_sig(1969)	<=	CN_out_sig(1619);
VN_in_sig(3021)	<=	CN_out_sig(1620);
VN_in_sig(3509)	<=	CN_out_sig(1621);
VN_in_sig(4065)	<=	CN_out_sig(1622);
VN_in_sig(5021)	<=	CN_out_sig(1623);
VN_in_sig(57)	<=	CN_out_sig(1624);
VN_in_sig(949)	<=	CN_out_sig(1625);
VN_in_sig(1325)	<=	CN_out_sig(1626);
VN_in_sig(1973)	<=	CN_out_sig(1627);
VN_in_sig(2809)	<=	CN_out_sig(1628);
VN_in_sig(3513)	<=	CN_out_sig(1629);
VN_in_sig(4069)	<=	CN_out_sig(1630);
VN_in_sig(5025)	<=	CN_out_sig(1631);
VN_in_sig(61)	<=	CN_out_sig(1632);
VN_in_sig(953)	<=	CN_out_sig(1633);
VN_in_sig(1329)	<=	CN_out_sig(1634);
VN_in_sig(1977)	<=	CN_out_sig(1635);
VN_in_sig(2813)	<=	CN_out_sig(1636);
VN_in_sig(3517)	<=	CN_out_sig(1637);
VN_in_sig(4073)	<=	CN_out_sig(1638);
VN_in_sig(5029)	<=	CN_out_sig(1639);
VN_in_sig(65)	<=	CN_out_sig(1640);
VN_in_sig(957)	<=	CN_out_sig(1641);
VN_in_sig(1333)	<=	CN_out_sig(1642);
VN_in_sig(1981)	<=	CN_out_sig(1643);
VN_in_sig(2817)	<=	CN_out_sig(1644);
VN_in_sig(3521)	<=	CN_out_sig(1645);
VN_in_sig(4077)	<=	CN_out_sig(1646);
VN_in_sig(5033)	<=	CN_out_sig(1647);
VN_in_sig(69)	<=	CN_out_sig(1648);
VN_in_sig(961)	<=	CN_out_sig(1649);
VN_in_sig(1337)	<=	CN_out_sig(1650);
VN_in_sig(1985)	<=	CN_out_sig(1651);
VN_in_sig(2821)	<=	CN_out_sig(1652);
VN_in_sig(3525)	<=	CN_out_sig(1653);
VN_in_sig(4081)	<=	CN_out_sig(1654);
VN_in_sig(5037)	<=	CN_out_sig(1655);
VN_in_sig(73)	<=	CN_out_sig(1656);
VN_in_sig(965)	<=	CN_out_sig(1657);
VN_in_sig(1341)	<=	CN_out_sig(1658);
VN_in_sig(1989)	<=	CN_out_sig(1659);
VN_in_sig(2825)	<=	CN_out_sig(1660);
VN_in_sig(3529)	<=	CN_out_sig(1661);
VN_in_sig(4085)	<=	CN_out_sig(1662);
VN_in_sig(5041)	<=	CN_out_sig(1663);
VN_in_sig(77)	<=	CN_out_sig(1664);
VN_in_sig(969)	<=	CN_out_sig(1665);
VN_in_sig(1345)	<=	CN_out_sig(1666);
VN_in_sig(1993)	<=	CN_out_sig(1667);
VN_in_sig(2829)	<=	CN_out_sig(1668);
VN_in_sig(3533)	<=	CN_out_sig(1669);
VN_in_sig(4089)	<=	CN_out_sig(1670);
VN_in_sig(5045)	<=	CN_out_sig(1671);
VN_in_sig(81)	<=	CN_out_sig(1672);
VN_in_sig(973)	<=	CN_out_sig(1673);
VN_in_sig(1349)	<=	CN_out_sig(1674);
VN_in_sig(1997)	<=	CN_out_sig(1675);
VN_in_sig(2833)	<=	CN_out_sig(1676);
VN_in_sig(3537)	<=	CN_out_sig(1677);
VN_in_sig(4093)	<=	CN_out_sig(1678);
VN_in_sig(5049)	<=	CN_out_sig(1679);
VN_in_sig(85)	<=	CN_out_sig(1680);
VN_in_sig(977)	<=	CN_out_sig(1681);
VN_in_sig(1353)	<=	CN_out_sig(1682);
VN_in_sig(2001)	<=	CN_out_sig(1683);
VN_in_sig(2837)	<=	CN_out_sig(1684);
VN_in_sig(3541)	<=	CN_out_sig(1685);
VN_in_sig(4097)	<=	CN_out_sig(1686);
VN_in_sig(5053)	<=	CN_out_sig(1687);
VN_in_sig(89)	<=	CN_out_sig(1688);
VN_in_sig(981)	<=	CN_out_sig(1689);
VN_in_sig(1357)	<=	CN_out_sig(1690);
VN_in_sig(2005)	<=	CN_out_sig(1691);
VN_in_sig(2841)	<=	CN_out_sig(1692);
VN_in_sig(3545)	<=	CN_out_sig(1693);
VN_in_sig(4101)	<=	CN_out_sig(1694);
VN_in_sig(5057)	<=	CN_out_sig(1695);
VN_in_sig(93)	<=	CN_out_sig(1696);
VN_in_sig(985)	<=	CN_out_sig(1697);
VN_in_sig(1361)	<=	CN_out_sig(1698);
VN_in_sig(2009)	<=	CN_out_sig(1699);
VN_in_sig(2845)	<=	CN_out_sig(1700);
VN_in_sig(3549)	<=	CN_out_sig(1701);
VN_in_sig(3889)	<=	CN_out_sig(1702);
VN_in_sig(5061)	<=	CN_out_sig(1703);
VN_in_sig(97)	<=	CN_out_sig(1704);
VN_in_sig(989)	<=	CN_out_sig(1705);
VN_in_sig(1365)	<=	CN_out_sig(1706);
VN_in_sig(2013)	<=	CN_out_sig(1707);
VN_in_sig(2849)	<=	CN_out_sig(1708);
VN_in_sig(3553)	<=	CN_out_sig(1709);
VN_in_sig(3893)	<=	CN_out_sig(1710);
VN_in_sig(5065)	<=	CN_out_sig(1711);
VN_in_sig(101)	<=	CN_out_sig(1712);
VN_in_sig(993)	<=	CN_out_sig(1713);
VN_in_sig(1369)	<=	CN_out_sig(1714);
VN_in_sig(2017)	<=	CN_out_sig(1715);
VN_in_sig(2853)	<=	CN_out_sig(1716);
VN_in_sig(3557)	<=	CN_out_sig(1717);
VN_in_sig(3897)	<=	CN_out_sig(1718);
VN_in_sig(5069)	<=	CN_out_sig(1719);
VN_in_sig(105)	<=	CN_out_sig(1720);
VN_in_sig(997)	<=	CN_out_sig(1721);
VN_in_sig(1373)	<=	CN_out_sig(1722);
VN_in_sig(2021)	<=	CN_out_sig(1723);
VN_in_sig(2857)	<=	CN_out_sig(1724);
VN_in_sig(3561)	<=	CN_out_sig(1725);
VN_in_sig(3901)	<=	CN_out_sig(1726);
VN_in_sig(5073)	<=	CN_out_sig(1727);
VN_in_sig(385)	<=	CN_out_sig(1728);
VN_in_sig(737)	<=	CN_out_sig(1729);
VN_in_sig(1557)	<=	CN_out_sig(1730);
VN_in_sig(2553)	<=	CN_out_sig(1731);
VN_in_sig(3041)	<=	CN_out_sig(1732);
VN_in_sig(3297)	<=	CN_out_sig(1733);
VN_in_sig(4501)	<=	CN_out_sig(1734);
VN_in_sig(4605)	<=	CN_out_sig(1735);
VN_in_sig(389)	<=	CN_out_sig(1736);
VN_in_sig(741)	<=	CN_out_sig(1737);
VN_in_sig(1561)	<=	CN_out_sig(1738);
VN_in_sig(2557)	<=	CN_out_sig(1739);
VN_in_sig(3045)	<=	CN_out_sig(1740);
VN_in_sig(3301)	<=	CN_out_sig(1741);
VN_in_sig(4505)	<=	CN_out_sig(1742);
VN_in_sig(4609)	<=	CN_out_sig(1743);
VN_in_sig(393)	<=	CN_out_sig(1744);
VN_in_sig(745)	<=	CN_out_sig(1745);
VN_in_sig(1565)	<=	CN_out_sig(1746);
VN_in_sig(2561)	<=	CN_out_sig(1747);
VN_in_sig(3049)	<=	CN_out_sig(1748);
VN_in_sig(3305)	<=	CN_out_sig(1749);
VN_in_sig(4509)	<=	CN_out_sig(1750);
VN_in_sig(4613)	<=	CN_out_sig(1751);
VN_in_sig(397)	<=	CN_out_sig(1752);
VN_in_sig(749)	<=	CN_out_sig(1753);
VN_in_sig(1569)	<=	CN_out_sig(1754);
VN_in_sig(2565)	<=	CN_out_sig(1755);
VN_in_sig(3053)	<=	CN_out_sig(1756);
VN_in_sig(3309)	<=	CN_out_sig(1757);
VN_in_sig(4513)	<=	CN_out_sig(1758);
VN_in_sig(4617)	<=	CN_out_sig(1759);
VN_in_sig(401)	<=	CN_out_sig(1760);
VN_in_sig(753)	<=	CN_out_sig(1761);
VN_in_sig(1573)	<=	CN_out_sig(1762);
VN_in_sig(2569)	<=	CN_out_sig(1763);
VN_in_sig(3057)	<=	CN_out_sig(1764);
VN_in_sig(3313)	<=	CN_out_sig(1765);
VN_in_sig(4517)	<=	CN_out_sig(1766);
VN_in_sig(4621)	<=	CN_out_sig(1767);
VN_in_sig(405)	<=	CN_out_sig(1768);
VN_in_sig(757)	<=	CN_out_sig(1769);
VN_in_sig(1577)	<=	CN_out_sig(1770);
VN_in_sig(2573)	<=	CN_out_sig(1771);
VN_in_sig(3061)	<=	CN_out_sig(1772);
VN_in_sig(3317)	<=	CN_out_sig(1773);
VN_in_sig(4521)	<=	CN_out_sig(1774);
VN_in_sig(4625)	<=	CN_out_sig(1775);
VN_in_sig(409)	<=	CN_out_sig(1776);
VN_in_sig(761)	<=	CN_out_sig(1777);
VN_in_sig(1581)	<=	CN_out_sig(1778);
VN_in_sig(2577)	<=	CN_out_sig(1779);
VN_in_sig(3065)	<=	CN_out_sig(1780);
VN_in_sig(3321)	<=	CN_out_sig(1781);
VN_in_sig(4525)	<=	CN_out_sig(1782);
VN_in_sig(4629)	<=	CN_out_sig(1783);
VN_in_sig(413)	<=	CN_out_sig(1784);
VN_in_sig(765)	<=	CN_out_sig(1785);
VN_in_sig(1585)	<=	CN_out_sig(1786);
VN_in_sig(2581)	<=	CN_out_sig(1787);
VN_in_sig(3069)	<=	CN_out_sig(1788);
VN_in_sig(3325)	<=	CN_out_sig(1789);
VN_in_sig(4529)	<=	CN_out_sig(1790);
VN_in_sig(4633)	<=	CN_out_sig(1791);
VN_in_sig(417)	<=	CN_out_sig(1792);
VN_in_sig(769)	<=	CN_out_sig(1793);
VN_in_sig(1589)	<=	CN_out_sig(1794);
VN_in_sig(2585)	<=	CN_out_sig(1795);
VN_in_sig(3073)	<=	CN_out_sig(1796);
VN_in_sig(3329)	<=	CN_out_sig(1797);
VN_in_sig(4533)	<=	CN_out_sig(1798);
VN_in_sig(4637)	<=	CN_out_sig(1799);
VN_in_sig(421)	<=	CN_out_sig(1800);
VN_in_sig(773)	<=	CN_out_sig(1801);
VN_in_sig(1593)	<=	CN_out_sig(1802);
VN_in_sig(2589)	<=	CN_out_sig(1803);
VN_in_sig(3077)	<=	CN_out_sig(1804);
VN_in_sig(3333)	<=	CN_out_sig(1805);
VN_in_sig(4321)	<=	CN_out_sig(1806);
VN_in_sig(4641)	<=	CN_out_sig(1807);
VN_in_sig(425)	<=	CN_out_sig(1808);
VN_in_sig(777)	<=	CN_out_sig(1809);
VN_in_sig(1597)	<=	CN_out_sig(1810);
VN_in_sig(2377)	<=	CN_out_sig(1811);
VN_in_sig(3081)	<=	CN_out_sig(1812);
VN_in_sig(3337)	<=	CN_out_sig(1813);
VN_in_sig(4325)	<=	CN_out_sig(1814);
VN_in_sig(4645)	<=	CN_out_sig(1815);
VN_in_sig(429)	<=	CN_out_sig(1816);
VN_in_sig(781)	<=	CN_out_sig(1817);
VN_in_sig(1601)	<=	CN_out_sig(1818);
VN_in_sig(2381)	<=	CN_out_sig(1819);
VN_in_sig(3085)	<=	CN_out_sig(1820);
VN_in_sig(3341)	<=	CN_out_sig(1821);
VN_in_sig(4329)	<=	CN_out_sig(1822);
VN_in_sig(4649)	<=	CN_out_sig(1823);
VN_in_sig(217)	<=	CN_out_sig(1824);
VN_in_sig(785)	<=	CN_out_sig(1825);
VN_in_sig(1605)	<=	CN_out_sig(1826);
VN_in_sig(2385)	<=	CN_out_sig(1827);
VN_in_sig(3089)	<=	CN_out_sig(1828);
VN_in_sig(3345)	<=	CN_out_sig(1829);
VN_in_sig(4333)	<=	CN_out_sig(1830);
VN_in_sig(4653)	<=	CN_out_sig(1831);
VN_in_sig(221)	<=	CN_out_sig(1832);
VN_in_sig(789)	<=	CN_out_sig(1833);
VN_in_sig(1609)	<=	CN_out_sig(1834);
VN_in_sig(2389)	<=	CN_out_sig(1835);
VN_in_sig(3093)	<=	CN_out_sig(1836);
VN_in_sig(3349)	<=	CN_out_sig(1837);
VN_in_sig(4337)	<=	CN_out_sig(1838);
VN_in_sig(4657)	<=	CN_out_sig(1839);
VN_in_sig(225)	<=	CN_out_sig(1840);
VN_in_sig(793)	<=	CN_out_sig(1841);
VN_in_sig(1613)	<=	CN_out_sig(1842);
VN_in_sig(2393)	<=	CN_out_sig(1843);
VN_in_sig(3097)	<=	CN_out_sig(1844);
VN_in_sig(3353)	<=	CN_out_sig(1845);
VN_in_sig(4341)	<=	CN_out_sig(1846);
VN_in_sig(4661)	<=	CN_out_sig(1847);
VN_in_sig(229)	<=	CN_out_sig(1848);
VN_in_sig(797)	<=	CN_out_sig(1849);
VN_in_sig(1617)	<=	CN_out_sig(1850);
VN_in_sig(2397)	<=	CN_out_sig(1851);
VN_in_sig(3101)	<=	CN_out_sig(1852);
VN_in_sig(3357)	<=	CN_out_sig(1853);
VN_in_sig(4345)	<=	CN_out_sig(1854);
VN_in_sig(4665)	<=	CN_out_sig(1855);
VN_in_sig(233)	<=	CN_out_sig(1856);
VN_in_sig(801)	<=	CN_out_sig(1857);
VN_in_sig(1621)	<=	CN_out_sig(1858);
VN_in_sig(2401)	<=	CN_out_sig(1859);
VN_in_sig(3105)	<=	CN_out_sig(1860);
VN_in_sig(3361)	<=	CN_out_sig(1861);
VN_in_sig(4349)	<=	CN_out_sig(1862);
VN_in_sig(4669)	<=	CN_out_sig(1863);
VN_in_sig(237)	<=	CN_out_sig(1864);
VN_in_sig(805)	<=	CN_out_sig(1865);
VN_in_sig(1625)	<=	CN_out_sig(1866);
VN_in_sig(2405)	<=	CN_out_sig(1867);
VN_in_sig(3109)	<=	CN_out_sig(1868);
VN_in_sig(3365)	<=	CN_out_sig(1869);
VN_in_sig(4353)	<=	CN_out_sig(1870);
VN_in_sig(4673)	<=	CN_out_sig(1871);
VN_in_sig(241)	<=	CN_out_sig(1872);
VN_in_sig(809)	<=	CN_out_sig(1873);
VN_in_sig(1629)	<=	CN_out_sig(1874);
VN_in_sig(2409)	<=	CN_out_sig(1875);
VN_in_sig(3113)	<=	CN_out_sig(1876);
VN_in_sig(3369)	<=	CN_out_sig(1877);
VN_in_sig(4357)	<=	CN_out_sig(1878);
VN_in_sig(4677)	<=	CN_out_sig(1879);
VN_in_sig(245)	<=	CN_out_sig(1880);
VN_in_sig(813)	<=	CN_out_sig(1881);
VN_in_sig(1633)	<=	CN_out_sig(1882);
VN_in_sig(2413)	<=	CN_out_sig(1883);
VN_in_sig(3117)	<=	CN_out_sig(1884);
VN_in_sig(3373)	<=	CN_out_sig(1885);
VN_in_sig(4361)	<=	CN_out_sig(1886);
VN_in_sig(4681)	<=	CN_out_sig(1887);
VN_in_sig(249)	<=	CN_out_sig(1888);
VN_in_sig(817)	<=	CN_out_sig(1889);
VN_in_sig(1637)	<=	CN_out_sig(1890);
VN_in_sig(2417)	<=	CN_out_sig(1891);
VN_in_sig(3121)	<=	CN_out_sig(1892);
VN_in_sig(3377)	<=	CN_out_sig(1893);
VN_in_sig(4365)	<=	CN_out_sig(1894);
VN_in_sig(4685)	<=	CN_out_sig(1895);
VN_in_sig(253)	<=	CN_out_sig(1896);
VN_in_sig(821)	<=	CN_out_sig(1897);
VN_in_sig(1641)	<=	CN_out_sig(1898);
VN_in_sig(2421)	<=	CN_out_sig(1899);
VN_in_sig(3125)	<=	CN_out_sig(1900);
VN_in_sig(3381)	<=	CN_out_sig(1901);
VN_in_sig(4369)	<=	CN_out_sig(1902);
VN_in_sig(4689)	<=	CN_out_sig(1903);
VN_in_sig(257)	<=	CN_out_sig(1904);
VN_in_sig(825)	<=	CN_out_sig(1905);
VN_in_sig(1645)	<=	CN_out_sig(1906);
VN_in_sig(2425)	<=	CN_out_sig(1907);
VN_in_sig(3129)	<=	CN_out_sig(1908);
VN_in_sig(3385)	<=	CN_out_sig(1909);
VN_in_sig(4373)	<=	CN_out_sig(1910);
VN_in_sig(4693)	<=	CN_out_sig(1911);
VN_in_sig(261)	<=	CN_out_sig(1912);
VN_in_sig(829)	<=	CN_out_sig(1913);
VN_in_sig(1649)	<=	CN_out_sig(1914);
VN_in_sig(2429)	<=	CN_out_sig(1915);
VN_in_sig(3133)	<=	CN_out_sig(1916);
VN_in_sig(3389)	<=	CN_out_sig(1917);
VN_in_sig(4377)	<=	CN_out_sig(1918);
VN_in_sig(4697)	<=	CN_out_sig(1919);
VN_in_sig(265)	<=	CN_out_sig(1920);
VN_in_sig(833)	<=	CN_out_sig(1921);
VN_in_sig(1653)	<=	CN_out_sig(1922);
VN_in_sig(2433)	<=	CN_out_sig(1923);
VN_in_sig(3137)	<=	CN_out_sig(1924);
VN_in_sig(3393)	<=	CN_out_sig(1925);
VN_in_sig(4381)	<=	CN_out_sig(1926);
VN_in_sig(4701)	<=	CN_out_sig(1927);
VN_in_sig(269)	<=	CN_out_sig(1928);
VN_in_sig(837)	<=	CN_out_sig(1929);
VN_in_sig(1657)	<=	CN_out_sig(1930);
VN_in_sig(2437)	<=	CN_out_sig(1931);
VN_in_sig(3141)	<=	CN_out_sig(1932);
VN_in_sig(3397)	<=	CN_out_sig(1933);
VN_in_sig(4385)	<=	CN_out_sig(1934);
VN_in_sig(4705)	<=	CN_out_sig(1935);
VN_in_sig(273)	<=	CN_out_sig(1936);
VN_in_sig(841)	<=	CN_out_sig(1937);
VN_in_sig(1661)	<=	CN_out_sig(1938);
VN_in_sig(2441)	<=	CN_out_sig(1939);
VN_in_sig(3145)	<=	CN_out_sig(1940);
VN_in_sig(3401)	<=	CN_out_sig(1941);
VN_in_sig(4389)	<=	CN_out_sig(1942);
VN_in_sig(4709)	<=	CN_out_sig(1943);
VN_in_sig(277)	<=	CN_out_sig(1944);
VN_in_sig(845)	<=	CN_out_sig(1945);
VN_in_sig(1665)	<=	CN_out_sig(1946);
VN_in_sig(2445)	<=	CN_out_sig(1947);
VN_in_sig(3149)	<=	CN_out_sig(1948);
VN_in_sig(3405)	<=	CN_out_sig(1949);
VN_in_sig(4393)	<=	CN_out_sig(1950);
VN_in_sig(4713)	<=	CN_out_sig(1951);
VN_in_sig(281)	<=	CN_out_sig(1952);
VN_in_sig(849)	<=	CN_out_sig(1953);
VN_in_sig(1669)	<=	CN_out_sig(1954);
VN_in_sig(2449)	<=	CN_out_sig(1955);
VN_in_sig(3153)	<=	CN_out_sig(1956);
VN_in_sig(3409)	<=	CN_out_sig(1957);
VN_in_sig(4397)	<=	CN_out_sig(1958);
VN_in_sig(4717)	<=	CN_out_sig(1959);
VN_in_sig(285)	<=	CN_out_sig(1960);
VN_in_sig(853)	<=	CN_out_sig(1961);
VN_in_sig(1673)	<=	CN_out_sig(1962);
VN_in_sig(2453)	<=	CN_out_sig(1963);
VN_in_sig(3157)	<=	CN_out_sig(1964);
VN_in_sig(3413)	<=	CN_out_sig(1965);
VN_in_sig(4401)	<=	CN_out_sig(1966);
VN_in_sig(4721)	<=	CN_out_sig(1967);
VN_in_sig(289)	<=	CN_out_sig(1968);
VN_in_sig(857)	<=	CN_out_sig(1969);
VN_in_sig(1677)	<=	CN_out_sig(1970);
VN_in_sig(2457)	<=	CN_out_sig(1971);
VN_in_sig(3161)	<=	CN_out_sig(1972);
VN_in_sig(3417)	<=	CN_out_sig(1973);
VN_in_sig(4405)	<=	CN_out_sig(1974);
VN_in_sig(4725)	<=	CN_out_sig(1975);
VN_in_sig(293)	<=	CN_out_sig(1976);
VN_in_sig(861)	<=	CN_out_sig(1977);
VN_in_sig(1681)	<=	CN_out_sig(1978);
VN_in_sig(2461)	<=	CN_out_sig(1979);
VN_in_sig(3165)	<=	CN_out_sig(1980);
VN_in_sig(3421)	<=	CN_out_sig(1981);
VN_in_sig(4409)	<=	CN_out_sig(1982);
VN_in_sig(4729)	<=	CN_out_sig(1983);
VN_in_sig(297)	<=	CN_out_sig(1984);
VN_in_sig(649)	<=	CN_out_sig(1985);
VN_in_sig(1685)	<=	CN_out_sig(1986);
VN_in_sig(2465)	<=	CN_out_sig(1987);
VN_in_sig(3169)	<=	CN_out_sig(1988);
VN_in_sig(3425)	<=	CN_out_sig(1989);
VN_in_sig(4413)	<=	CN_out_sig(1990);
VN_in_sig(4733)	<=	CN_out_sig(1991);
VN_in_sig(301)	<=	CN_out_sig(1992);
VN_in_sig(653)	<=	CN_out_sig(1993);
VN_in_sig(1689)	<=	CN_out_sig(1994);
VN_in_sig(2469)	<=	CN_out_sig(1995);
VN_in_sig(3173)	<=	CN_out_sig(1996);
VN_in_sig(3429)	<=	CN_out_sig(1997);
VN_in_sig(4417)	<=	CN_out_sig(1998);
VN_in_sig(4737)	<=	CN_out_sig(1999);
VN_in_sig(305)	<=	CN_out_sig(2000);
VN_in_sig(657)	<=	CN_out_sig(2001);
VN_in_sig(1693)	<=	CN_out_sig(2002);
VN_in_sig(2473)	<=	CN_out_sig(2003);
VN_in_sig(3177)	<=	CN_out_sig(2004);
VN_in_sig(3433)	<=	CN_out_sig(2005);
VN_in_sig(4421)	<=	CN_out_sig(2006);
VN_in_sig(4741)	<=	CN_out_sig(2007);
VN_in_sig(309)	<=	CN_out_sig(2008);
VN_in_sig(661)	<=	CN_out_sig(2009);
VN_in_sig(1697)	<=	CN_out_sig(2010);
VN_in_sig(2477)	<=	CN_out_sig(2011);
VN_in_sig(3181)	<=	CN_out_sig(2012);
VN_in_sig(3437)	<=	CN_out_sig(2013);
VN_in_sig(4425)	<=	CN_out_sig(2014);
VN_in_sig(4745)	<=	CN_out_sig(2015);
VN_in_sig(313)	<=	CN_out_sig(2016);
VN_in_sig(665)	<=	CN_out_sig(2017);
VN_in_sig(1701)	<=	CN_out_sig(2018);
VN_in_sig(2481)	<=	CN_out_sig(2019);
VN_in_sig(3185)	<=	CN_out_sig(2020);
VN_in_sig(3441)	<=	CN_out_sig(2021);
VN_in_sig(4429)	<=	CN_out_sig(2022);
VN_in_sig(4749)	<=	CN_out_sig(2023);
VN_in_sig(317)	<=	CN_out_sig(2024);
VN_in_sig(669)	<=	CN_out_sig(2025);
VN_in_sig(1705)	<=	CN_out_sig(2026);
VN_in_sig(2485)	<=	CN_out_sig(2027);
VN_in_sig(3189)	<=	CN_out_sig(2028);
VN_in_sig(3445)	<=	CN_out_sig(2029);
VN_in_sig(4433)	<=	CN_out_sig(2030);
VN_in_sig(4537)	<=	CN_out_sig(2031);
VN_in_sig(321)	<=	CN_out_sig(2032);
VN_in_sig(673)	<=	CN_out_sig(2033);
VN_in_sig(1709)	<=	CN_out_sig(2034);
VN_in_sig(2489)	<=	CN_out_sig(2035);
VN_in_sig(3193)	<=	CN_out_sig(2036);
VN_in_sig(3449)	<=	CN_out_sig(2037);
VN_in_sig(4437)	<=	CN_out_sig(2038);
VN_in_sig(4541)	<=	CN_out_sig(2039);
VN_in_sig(325)	<=	CN_out_sig(2040);
VN_in_sig(677)	<=	CN_out_sig(2041);
VN_in_sig(1713)	<=	CN_out_sig(2042);
VN_in_sig(2493)	<=	CN_out_sig(2043);
VN_in_sig(3197)	<=	CN_out_sig(2044);
VN_in_sig(3453)	<=	CN_out_sig(2045);
VN_in_sig(4441)	<=	CN_out_sig(2046);
VN_in_sig(4545)	<=	CN_out_sig(2047);
VN_in_sig(329)	<=	CN_out_sig(2048);
VN_in_sig(681)	<=	CN_out_sig(2049);
VN_in_sig(1717)	<=	CN_out_sig(2050);
VN_in_sig(2497)	<=	CN_out_sig(2051);
VN_in_sig(3201)	<=	CN_out_sig(2052);
VN_in_sig(3241)	<=	CN_out_sig(2053);
VN_in_sig(4445)	<=	CN_out_sig(2054);
VN_in_sig(4549)	<=	CN_out_sig(2055);
VN_in_sig(333)	<=	CN_out_sig(2056);
VN_in_sig(685)	<=	CN_out_sig(2057);
VN_in_sig(1721)	<=	CN_out_sig(2058);
VN_in_sig(2501)	<=	CN_out_sig(2059);
VN_in_sig(3205)	<=	CN_out_sig(2060);
VN_in_sig(3245)	<=	CN_out_sig(2061);
VN_in_sig(4449)	<=	CN_out_sig(2062);
VN_in_sig(4553)	<=	CN_out_sig(2063);
VN_in_sig(337)	<=	CN_out_sig(2064);
VN_in_sig(689)	<=	CN_out_sig(2065);
VN_in_sig(1725)	<=	CN_out_sig(2066);
VN_in_sig(2505)	<=	CN_out_sig(2067);
VN_in_sig(3209)	<=	CN_out_sig(2068);
VN_in_sig(3249)	<=	CN_out_sig(2069);
VN_in_sig(4453)	<=	CN_out_sig(2070);
VN_in_sig(4557)	<=	CN_out_sig(2071);
VN_in_sig(341)	<=	CN_out_sig(2072);
VN_in_sig(693)	<=	CN_out_sig(2073);
VN_in_sig(1513)	<=	CN_out_sig(2074);
VN_in_sig(2509)	<=	CN_out_sig(2075);
VN_in_sig(3213)	<=	CN_out_sig(2076);
VN_in_sig(3253)	<=	CN_out_sig(2077);
VN_in_sig(4457)	<=	CN_out_sig(2078);
VN_in_sig(4561)	<=	CN_out_sig(2079);
VN_in_sig(345)	<=	CN_out_sig(2080);
VN_in_sig(697)	<=	CN_out_sig(2081);
VN_in_sig(1517)	<=	CN_out_sig(2082);
VN_in_sig(2513)	<=	CN_out_sig(2083);
VN_in_sig(3217)	<=	CN_out_sig(2084);
VN_in_sig(3257)	<=	CN_out_sig(2085);
VN_in_sig(4461)	<=	CN_out_sig(2086);
VN_in_sig(4565)	<=	CN_out_sig(2087);
VN_in_sig(349)	<=	CN_out_sig(2088);
VN_in_sig(701)	<=	CN_out_sig(2089);
VN_in_sig(1521)	<=	CN_out_sig(2090);
VN_in_sig(2517)	<=	CN_out_sig(2091);
VN_in_sig(3221)	<=	CN_out_sig(2092);
VN_in_sig(3261)	<=	CN_out_sig(2093);
VN_in_sig(4465)	<=	CN_out_sig(2094);
VN_in_sig(4569)	<=	CN_out_sig(2095);
VN_in_sig(353)	<=	CN_out_sig(2096);
VN_in_sig(705)	<=	CN_out_sig(2097);
VN_in_sig(1525)	<=	CN_out_sig(2098);
VN_in_sig(2521)	<=	CN_out_sig(2099);
VN_in_sig(3225)	<=	CN_out_sig(2100);
VN_in_sig(3265)	<=	CN_out_sig(2101);
VN_in_sig(4469)	<=	CN_out_sig(2102);
VN_in_sig(4573)	<=	CN_out_sig(2103);
VN_in_sig(357)	<=	CN_out_sig(2104);
VN_in_sig(709)	<=	CN_out_sig(2105);
VN_in_sig(1529)	<=	CN_out_sig(2106);
VN_in_sig(2525)	<=	CN_out_sig(2107);
VN_in_sig(3229)	<=	CN_out_sig(2108);
VN_in_sig(3269)	<=	CN_out_sig(2109);
VN_in_sig(4473)	<=	CN_out_sig(2110);
VN_in_sig(4577)	<=	CN_out_sig(2111);
VN_in_sig(361)	<=	CN_out_sig(2112);
VN_in_sig(713)	<=	CN_out_sig(2113);
VN_in_sig(1533)	<=	CN_out_sig(2114);
VN_in_sig(2529)	<=	CN_out_sig(2115);
VN_in_sig(3233)	<=	CN_out_sig(2116);
VN_in_sig(3273)	<=	CN_out_sig(2117);
VN_in_sig(4477)	<=	CN_out_sig(2118);
VN_in_sig(4581)	<=	CN_out_sig(2119);
VN_in_sig(365)	<=	CN_out_sig(2120);
VN_in_sig(717)	<=	CN_out_sig(2121);
VN_in_sig(1537)	<=	CN_out_sig(2122);
VN_in_sig(2533)	<=	CN_out_sig(2123);
VN_in_sig(3237)	<=	CN_out_sig(2124);
VN_in_sig(3277)	<=	CN_out_sig(2125);
VN_in_sig(4481)	<=	CN_out_sig(2126);
VN_in_sig(4585)	<=	CN_out_sig(2127);
VN_in_sig(369)	<=	CN_out_sig(2128);
VN_in_sig(721)	<=	CN_out_sig(2129);
VN_in_sig(1541)	<=	CN_out_sig(2130);
VN_in_sig(2537)	<=	CN_out_sig(2131);
VN_in_sig(3025)	<=	CN_out_sig(2132);
VN_in_sig(3281)	<=	CN_out_sig(2133);
VN_in_sig(4485)	<=	CN_out_sig(2134);
VN_in_sig(4589)	<=	CN_out_sig(2135);
VN_in_sig(373)	<=	CN_out_sig(2136);
VN_in_sig(725)	<=	CN_out_sig(2137);
VN_in_sig(1545)	<=	CN_out_sig(2138);
VN_in_sig(2541)	<=	CN_out_sig(2139);
VN_in_sig(3029)	<=	CN_out_sig(2140);
VN_in_sig(3285)	<=	CN_out_sig(2141);
VN_in_sig(4489)	<=	CN_out_sig(2142);
VN_in_sig(4593)	<=	CN_out_sig(2143);
VN_in_sig(377)	<=	CN_out_sig(2144);
VN_in_sig(729)	<=	CN_out_sig(2145);
VN_in_sig(1549)	<=	CN_out_sig(2146);
VN_in_sig(2545)	<=	CN_out_sig(2147);
VN_in_sig(3033)	<=	CN_out_sig(2148);
VN_in_sig(3289)	<=	CN_out_sig(2149);
VN_in_sig(4493)	<=	CN_out_sig(2150);
VN_in_sig(4597)	<=	CN_out_sig(2151);
VN_in_sig(381)	<=	CN_out_sig(2152);
VN_in_sig(733)	<=	CN_out_sig(2153);
VN_in_sig(1553)	<=	CN_out_sig(2154);
VN_in_sig(2549)	<=	CN_out_sig(2155);
VN_in_sig(3037)	<=	CN_out_sig(2156);
VN_in_sig(3293)	<=	CN_out_sig(2157);
VN_in_sig(4497)	<=	CN_out_sig(2158);
VN_in_sig(4601)	<=	CN_out_sig(2159);
VN_in_sig(529)	<=	CN_out_sig(2160);
VN_in_sig(1121)	<=	CN_out_sig(2161);
VN_in_sig(1769)	<=	CN_out_sig(2162);
VN_in_sig(2233)	<=	CN_out_sig(2163);
VN_in_sig(2601)	<=	CN_out_sig(2164);
VN_in_sig(3749)	<=	CN_out_sig(2165);
VN_in_sig(4257)	<=	CN_out_sig(2166);
VN_in_sig(4877)	<=	CN_out_sig(2167);
VN_in_sig(533)	<=	CN_out_sig(2168);
VN_in_sig(1125)	<=	CN_out_sig(2169);
VN_in_sig(1773)	<=	CN_out_sig(2170);
VN_in_sig(2237)	<=	CN_out_sig(2171);
VN_in_sig(2605)	<=	CN_out_sig(2172);
VN_in_sig(3753)	<=	CN_out_sig(2173);
VN_in_sig(4261)	<=	CN_out_sig(2174);
VN_in_sig(4881)	<=	CN_out_sig(2175);
VN_in_sig(537)	<=	CN_out_sig(2176);
VN_in_sig(1129)	<=	CN_out_sig(2177);
VN_in_sig(1777)	<=	CN_out_sig(2178);
VN_in_sig(2241)	<=	CN_out_sig(2179);
VN_in_sig(2609)	<=	CN_out_sig(2180);
VN_in_sig(3757)	<=	CN_out_sig(2181);
VN_in_sig(4265)	<=	CN_out_sig(2182);
VN_in_sig(4885)	<=	CN_out_sig(2183);
VN_in_sig(541)	<=	CN_out_sig(2184);
VN_in_sig(1133)	<=	CN_out_sig(2185);
VN_in_sig(1781)	<=	CN_out_sig(2186);
VN_in_sig(2245)	<=	CN_out_sig(2187);
VN_in_sig(2613)	<=	CN_out_sig(2188);
VN_in_sig(3761)	<=	CN_out_sig(2189);
VN_in_sig(4269)	<=	CN_out_sig(2190);
VN_in_sig(4889)	<=	CN_out_sig(2191);
VN_in_sig(545)	<=	CN_out_sig(2192);
VN_in_sig(1137)	<=	CN_out_sig(2193);
VN_in_sig(1785)	<=	CN_out_sig(2194);
VN_in_sig(2249)	<=	CN_out_sig(2195);
VN_in_sig(2617)	<=	CN_out_sig(2196);
VN_in_sig(3765)	<=	CN_out_sig(2197);
VN_in_sig(4273)	<=	CN_out_sig(2198);
VN_in_sig(4893)	<=	CN_out_sig(2199);
VN_in_sig(549)	<=	CN_out_sig(2200);
VN_in_sig(1141)	<=	CN_out_sig(2201);
VN_in_sig(1789)	<=	CN_out_sig(2202);
VN_in_sig(2253)	<=	CN_out_sig(2203);
VN_in_sig(2621)	<=	CN_out_sig(2204);
VN_in_sig(3769)	<=	CN_out_sig(2205);
VN_in_sig(4277)	<=	CN_out_sig(2206);
VN_in_sig(4897)	<=	CN_out_sig(2207);
VN_in_sig(553)	<=	CN_out_sig(2208);
VN_in_sig(1145)	<=	CN_out_sig(2209);
VN_in_sig(1793)	<=	CN_out_sig(2210);
VN_in_sig(2257)	<=	CN_out_sig(2211);
VN_in_sig(2625)	<=	CN_out_sig(2212);
VN_in_sig(3773)	<=	CN_out_sig(2213);
VN_in_sig(4281)	<=	CN_out_sig(2214);
VN_in_sig(4901)	<=	CN_out_sig(2215);
VN_in_sig(557)	<=	CN_out_sig(2216);
VN_in_sig(1149)	<=	CN_out_sig(2217);
VN_in_sig(1797)	<=	CN_out_sig(2218);
VN_in_sig(2261)	<=	CN_out_sig(2219);
VN_in_sig(2629)	<=	CN_out_sig(2220);
VN_in_sig(3777)	<=	CN_out_sig(2221);
VN_in_sig(4285)	<=	CN_out_sig(2222);
VN_in_sig(4905)	<=	CN_out_sig(2223);
VN_in_sig(561)	<=	CN_out_sig(2224);
VN_in_sig(1153)	<=	CN_out_sig(2225);
VN_in_sig(1801)	<=	CN_out_sig(2226);
VN_in_sig(2265)	<=	CN_out_sig(2227);
VN_in_sig(2633)	<=	CN_out_sig(2228);
VN_in_sig(3781)	<=	CN_out_sig(2229);
VN_in_sig(4289)	<=	CN_out_sig(2230);
VN_in_sig(4909)	<=	CN_out_sig(2231);
VN_in_sig(565)	<=	CN_out_sig(2232);
VN_in_sig(1157)	<=	CN_out_sig(2233);
VN_in_sig(1805)	<=	CN_out_sig(2234);
VN_in_sig(2269)	<=	CN_out_sig(2235);
VN_in_sig(2637)	<=	CN_out_sig(2236);
VN_in_sig(3785)	<=	CN_out_sig(2237);
VN_in_sig(4293)	<=	CN_out_sig(2238);
VN_in_sig(4913)	<=	CN_out_sig(2239);
VN_in_sig(569)	<=	CN_out_sig(2240);
VN_in_sig(1161)	<=	CN_out_sig(2241);
VN_in_sig(1809)	<=	CN_out_sig(2242);
VN_in_sig(2273)	<=	CN_out_sig(2243);
VN_in_sig(2641)	<=	CN_out_sig(2244);
VN_in_sig(3789)	<=	CN_out_sig(2245);
VN_in_sig(4297)	<=	CN_out_sig(2246);
VN_in_sig(4917)	<=	CN_out_sig(2247);
VN_in_sig(573)	<=	CN_out_sig(2248);
VN_in_sig(1165)	<=	CN_out_sig(2249);
VN_in_sig(1813)	<=	CN_out_sig(2250);
VN_in_sig(2277)	<=	CN_out_sig(2251);
VN_in_sig(2645)	<=	CN_out_sig(2252);
VN_in_sig(3793)	<=	CN_out_sig(2253);
VN_in_sig(4301)	<=	CN_out_sig(2254);
VN_in_sig(4921)	<=	CN_out_sig(2255);
VN_in_sig(577)	<=	CN_out_sig(2256);
VN_in_sig(1169)	<=	CN_out_sig(2257);
VN_in_sig(1817)	<=	CN_out_sig(2258);
VN_in_sig(2281)	<=	CN_out_sig(2259);
VN_in_sig(2649)	<=	CN_out_sig(2260);
VN_in_sig(3797)	<=	CN_out_sig(2261);
VN_in_sig(4305)	<=	CN_out_sig(2262);
VN_in_sig(4925)	<=	CN_out_sig(2263);
VN_in_sig(581)	<=	CN_out_sig(2264);
VN_in_sig(1173)	<=	CN_out_sig(2265);
VN_in_sig(1821)	<=	CN_out_sig(2266);
VN_in_sig(2285)	<=	CN_out_sig(2267);
VN_in_sig(2653)	<=	CN_out_sig(2268);
VN_in_sig(3801)	<=	CN_out_sig(2269);
VN_in_sig(4309)	<=	CN_out_sig(2270);
VN_in_sig(4929)	<=	CN_out_sig(2271);
VN_in_sig(585)	<=	CN_out_sig(2272);
VN_in_sig(1177)	<=	CN_out_sig(2273);
VN_in_sig(1825)	<=	CN_out_sig(2274);
VN_in_sig(2289)	<=	CN_out_sig(2275);
VN_in_sig(2657)	<=	CN_out_sig(2276);
VN_in_sig(3805)	<=	CN_out_sig(2277);
VN_in_sig(4313)	<=	CN_out_sig(2278);
VN_in_sig(4933)	<=	CN_out_sig(2279);
VN_in_sig(589)	<=	CN_out_sig(2280);
VN_in_sig(1181)	<=	CN_out_sig(2281);
VN_in_sig(1829)	<=	CN_out_sig(2282);
VN_in_sig(2293)	<=	CN_out_sig(2283);
VN_in_sig(2661)	<=	CN_out_sig(2284);
VN_in_sig(3809)	<=	CN_out_sig(2285);
VN_in_sig(4317)	<=	CN_out_sig(2286);
VN_in_sig(4937)	<=	CN_out_sig(2287);
VN_in_sig(593)	<=	CN_out_sig(2288);
VN_in_sig(1185)	<=	CN_out_sig(2289);
VN_in_sig(1833)	<=	CN_out_sig(2290);
VN_in_sig(2297)	<=	CN_out_sig(2291);
VN_in_sig(2665)	<=	CN_out_sig(2292);
VN_in_sig(3813)	<=	CN_out_sig(2293);
VN_in_sig(4105)	<=	CN_out_sig(2294);
VN_in_sig(4941)	<=	CN_out_sig(2295);
VN_in_sig(597)	<=	CN_out_sig(2296);
VN_in_sig(1189)	<=	CN_out_sig(2297);
VN_in_sig(1837)	<=	CN_out_sig(2298);
VN_in_sig(2301)	<=	CN_out_sig(2299);
VN_in_sig(2669)	<=	CN_out_sig(2300);
VN_in_sig(3817)	<=	CN_out_sig(2301);
VN_in_sig(4109)	<=	CN_out_sig(2302);
VN_in_sig(4945)	<=	CN_out_sig(2303);
VN_in_sig(601)	<=	CN_out_sig(2304);
VN_in_sig(1193)	<=	CN_out_sig(2305);
VN_in_sig(1841)	<=	CN_out_sig(2306);
VN_in_sig(2305)	<=	CN_out_sig(2307);
VN_in_sig(2673)	<=	CN_out_sig(2308);
VN_in_sig(3821)	<=	CN_out_sig(2309);
VN_in_sig(4113)	<=	CN_out_sig(2310);
VN_in_sig(4949)	<=	CN_out_sig(2311);
VN_in_sig(605)	<=	CN_out_sig(2312);
VN_in_sig(1197)	<=	CN_out_sig(2313);
VN_in_sig(1845)	<=	CN_out_sig(2314);
VN_in_sig(2309)	<=	CN_out_sig(2315);
VN_in_sig(2677)	<=	CN_out_sig(2316);
VN_in_sig(3825)	<=	CN_out_sig(2317);
VN_in_sig(4117)	<=	CN_out_sig(2318);
VN_in_sig(4953)	<=	CN_out_sig(2319);
VN_in_sig(609)	<=	CN_out_sig(2320);
VN_in_sig(1201)	<=	CN_out_sig(2321);
VN_in_sig(1849)	<=	CN_out_sig(2322);
VN_in_sig(2313)	<=	CN_out_sig(2323);
VN_in_sig(2681)	<=	CN_out_sig(2324);
VN_in_sig(3829)	<=	CN_out_sig(2325);
VN_in_sig(4121)	<=	CN_out_sig(2326);
VN_in_sig(4957)	<=	CN_out_sig(2327);
VN_in_sig(613)	<=	CN_out_sig(2328);
VN_in_sig(1205)	<=	CN_out_sig(2329);
VN_in_sig(1853)	<=	CN_out_sig(2330);
VN_in_sig(2317)	<=	CN_out_sig(2331);
VN_in_sig(2685)	<=	CN_out_sig(2332);
VN_in_sig(3833)	<=	CN_out_sig(2333);
VN_in_sig(4125)	<=	CN_out_sig(2334);
VN_in_sig(4961)	<=	CN_out_sig(2335);
VN_in_sig(617)	<=	CN_out_sig(2336);
VN_in_sig(1209)	<=	CN_out_sig(2337);
VN_in_sig(1857)	<=	CN_out_sig(2338);
VN_in_sig(2321)	<=	CN_out_sig(2339);
VN_in_sig(2689)	<=	CN_out_sig(2340);
VN_in_sig(3837)	<=	CN_out_sig(2341);
VN_in_sig(4129)	<=	CN_out_sig(2342);
VN_in_sig(4965)	<=	CN_out_sig(2343);
VN_in_sig(621)	<=	CN_out_sig(2344);
VN_in_sig(1213)	<=	CN_out_sig(2345);
VN_in_sig(1861)	<=	CN_out_sig(2346);
VN_in_sig(2325)	<=	CN_out_sig(2347);
VN_in_sig(2693)	<=	CN_out_sig(2348);
VN_in_sig(3841)	<=	CN_out_sig(2349);
VN_in_sig(4133)	<=	CN_out_sig(2350);
VN_in_sig(4753)	<=	CN_out_sig(2351);
VN_in_sig(625)	<=	CN_out_sig(2352);
VN_in_sig(1217)	<=	CN_out_sig(2353);
VN_in_sig(1865)	<=	CN_out_sig(2354);
VN_in_sig(2329)	<=	CN_out_sig(2355);
VN_in_sig(2697)	<=	CN_out_sig(2356);
VN_in_sig(3845)	<=	CN_out_sig(2357);
VN_in_sig(4137)	<=	CN_out_sig(2358);
VN_in_sig(4757)	<=	CN_out_sig(2359);
VN_in_sig(629)	<=	CN_out_sig(2360);
VN_in_sig(1221)	<=	CN_out_sig(2361);
VN_in_sig(1869)	<=	CN_out_sig(2362);
VN_in_sig(2333)	<=	CN_out_sig(2363);
VN_in_sig(2701)	<=	CN_out_sig(2364);
VN_in_sig(3849)	<=	CN_out_sig(2365);
VN_in_sig(4141)	<=	CN_out_sig(2366);
VN_in_sig(4761)	<=	CN_out_sig(2367);
VN_in_sig(633)	<=	CN_out_sig(2368);
VN_in_sig(1225)	<=	CN_out_sig(2369);
VN_in_sig(1873)	<=	CN_out_sig(2370);
VN_in_sig(2337)	<=	CN_out_sig(2371);
VN_in_sig(2705)	<=	CN_out_sig(2372);
VN_in_sig(3853)	<=	CN_out_sig(2373);
VN_in_sig(4145)	<=	CN_out_sig(2374);
VN_in_sig(4765)	<=	CN_out_sig(2375);
VN_in_sig(637)	<=	CN_out_sig(2376);
VN_in_sig(1229)	<=	CN_out_sig(2377);
VN_in_sig(1877)	<=	CN_out_sig(2378);
VN_in_sig(2341)	<=	CN_out_sig(2379);
VN_in_sig(2709)	<=	CN_out_sig(2380);
VN_in_sig(3857)	<=	CN_out_sig(2381);
VN_in_sig(4149)	<=	CN_out_sig(2382);
VN_in_sig(4769)	<=	CN_out_sig(2383);
VN_in_sig(641)	<=	CN_out_sig(2384);
VN_in_sig(1233)	<=	CN_out_sig(2385);
VN_in_sig(1881)	<=	CN_out_sig(2386);
VN_in_sig(2345)	<=	CN_out_sig(2387);
VN_in_sig(2713)	<=	CN_out_sig(2388);
VN_in_sig(3861)	<=	CN_out_sig(2389);
VN_in_sig(4153)	<=	CN_out_sig(2390);
VN_in_sig(4773)	<=	CN_out_sig(2391);
VN_in_sig(645)	<=	CN_out_sig(2392);
VN_in_sig(1237)	<=	CN_out_sig(2393);
VN_in_sig(1885)	<=	CN_out_sig(2394);
VN_in_sig(2349)	<=	CN_out_sig(2395);
VN_in_sig(2717)	<=	CN_out_sig(2396);
VN_in_sig(3865)	<=	CN_out_sig(2397);
VN_in_sig(4157)	<=	CN_out_sig(2398);
VN_in_sig(4777)	<=	CN_out_sig(2399);
VN_in_sig(433)	<=	CN_out_sig(2400);
VN_in_sig(1241)	<=	CN_out_sig(2401);
VN_in_sig(1889)	<=	CN_out_sig(2402);
VN_in_sig(2353)	<=	CN_out_sig(2403);
VN_in_sig(2721)	<=	CN_out_sig(2404);
VN_in_sig(3869)	<=	CN_out_sig(2405);
VN_in_sig(4161)	<=	CN_out_sig(2406);
VN_in_sig(4781)	<=	CN_out_sig(2407);
VN_in_sig(437)	<=	CN_out_sig(2408);
VN_in_sig(1245)	<=	CN_out_sig(2409);
VN_in_sig(1893)	<=	CN_out_sig(2410);
VN_in_sig(2357)	<=	CN_out_sig(2411);
VN_in_sig(2725)	<=	CN_out_sig(2412);
VN_in_sig(3873)	<=	CN_out_sig(2413);
VN_in_sig(4165)	<=	CN_out_sig(2414);
VN_in_sig(4785)	<=	CN_out_sig(2415);
VN_in_sig(441)	<=	CN_out_sig(2416);
VN_in_sig(1249)	<=	CN_out_sig(2417);
VN_in_sig(1897)	<=	CN_out_sig(2418);
VN_in_sig(2361)	<=	CN_out_sig(2419);
VN_in_sig(2729)	<=	CN_out_sig(2420);
VN_in_sig(3877)	<=	CN_out_sig(2421);
VN_in_sig(4169)	<=	CN_out_sig(2422);
VN_in_sig(4789)	<=	CN_out_sig(2423);
VN_in_sig(445)	<=	CN_out_sig(2424);
VN_in_sig(1253)	<=	CN_out_sig(2425);
VN_in_sig(1901)	<=	CN_out_sig(2426);
VN_in_sig(2365)	<=	CN_out_sig(2427);
VN_in_sig(2733)	<=	CN_out_sig(2428);
VN_in_sig(3881)	<=	CN_out_sig(2429);
VN_in_sig(4173)	<=	CN_out_sig(2430);
VN_in_sig(4793)	<=	CN_out_sig(2431);
VN_in_sig(449)	<=	CN_out_sig(2432);
VN_in_sig(1257)	<=	CN_out_sig(2433);
VN_in_sig(1905)	<=	CN_out_sig(2434);
VN_in_sig(2369)	<=	CN_out_sig(2435);
VN_in_sig(2737)	<=	CN_out_sig(2436);
VN_in_sig(3885)	<=	CN_out_sig(2437);
VN_in_sig(4177)	<=	CN_out_sig(2438);
VN_in_sig(4797)	<=	CN_out_sig(2439);
VN_in_sig(453)	<=	CN_out_sig(2440);
VN_in_sig(1261)	<=	CN_out_sig(2441);
VN_in_sig(1909)	<=	CN_out_sig(2442);
VN_in_sig(2373)	<=	CN_out_sig(2443);
VN_in_sig(2741)	<=	CN_out_sig(2444);
VN_in_sig(3673)	<=	CN_out_sig(2445);
VN_in_sig(4181)	<=	CN_out_sig(2446);
VN_in_sig(4801)	<=	CN_out_sig(2447);
VN_in_sig(457)	<=	CN_out_sig(2448);
VN_in_sig(1265)	<=	CN_out_sig(2449);
VN_in_sig(1913)	<=	CN_out_sig(2450);
VN_in_sig(2161)	<=	CN_out_sig(2451);
VN_in_sig(2745)	<=	CN_out_sig(2452);
VN_in_sig(3677)	<=	CN_out_sig(2453);
VN_in_sig(4185)	<=	CN_out_sig(2454);
VN_in_sig(4805)	<=	CN_out_sig(2455);
VN_in_sig(461)	<=	CN_out_sig(2456);
VN_in_sig(1269)	<=	CN_out_sig(2457);
VN_in_sig(1917)	<=	CN_out_sig(2458);
VN_in_sig(2165)	<=	CN_out_sig(2459);
VN_in_sig(2749)	<=	CN_out_sig(2460);
VN_in_sig(3681)	<=	CN_out_sig(2461);
VN_in_sig(4189)	<=	CN_out_sig(2462);
VN_in_sig(4809)	<=	CN_out_sig(2463);
VN_in_sig(465)	<=	CN_out_sig(2464);
VN_in_sig(1273)	<=	CN_out_sig(2465);
VN_in_sig(1921)	<=	CN_out_sig(2466);
VN_in_sig(2169)	<=	CN_out_sig(2467);
VN_in_sig(2753)	<=	CN_out_sig(2468);
VN_in_sig(3685)	<=	CN_out_sig(2469);
VN_in_sig(4193)	<=	CN_out_sig(2470);
VN_in_sig(4813)	<=	CN_out_sig(2471);
VN_in_sig(469)	<=	CN_out_sig(2472);
VN_in_sig(1277)	<=	CN_out_sig(2473);
VN_in_sig(1925)	<=	CN_out_sig(2474);
VN_in_sig(2173)	<=	CN_out_sig(2475);
VN_in_sig(2757)	<=	CN_out_sig(2476);
VN_in_sig(3689)	<=	CN_out_sig(2477);
VN_in_sig(4197)	<=	CN_out_sig(2478);
VN_in_sig(4817)	<=	CN_out_sig(2479);
VN_in_sig(473)	<=	CN_out_sig(2480);
VN_in_sig(1281)	<=	CN_out_sig(2481);
VN_in_sig(1929)	<=	CN_out_sig(2482);
VN_in_sig(2177)	<=	CN_out_sig(2483);
VN_in_sig(2761)	<=	CN_out_sig(2484);
VN_in_sig(3693)	<=	CN_out_sig(2485);
VN_in_sig(4201)	<=	CN_out_sig(2486);
VN_in_sig(4821)	<=	CN_out_sig(2487);
VN_in_sig(477)	<=	CN_out_sig(2488);
VN_in_sig(1285)	<=	CN_out_sig(2489);
VN_in_sig(1933)	<=	CN_out_sig(2490);
VN_in_sig(2181)	<=	CN_out_sig(2491);
VN_in_sig(2765)	<=	CN_out_sig(2492);
VN_in_sig(3697)	<=	CN_out_sig(2493);
VN_in_sig(4205)	<=	CN_out_sig(2494);
VN_in_sig(4825)	<=	CN_out_sig(2495);
VN_in_sig(481)	<=	CN_out_sig(2496);
VN_in_sig(1289)	<=	CN_out_sig(2497);
VN_in_sig(1937)	<=	CN_out_sig(2498);
VN_in_sig(2185)	<=	CN_out_sig(2499);
VN_in_sig(2769)	<=	CN_out_sig(2500);
VN_in_sig(3701)	<=	CN_out_sig(2501);
VN_in_sig(4209)	<=	CN_out_sig(2502);
VN_in_sig(4829)	<=	CN_out_sig(2503);
VN_in_sig(485)	<=	CN_out_sig(2504);
VN_in_sig(1293)	<=	CN_out_sig(2505);
VN_in_sig(1941)	<=	CN_out_sig(2506);
VN_in_sig(2189)	<=	CN_out_sig(2507);
VN_in_sig(2773)	<=	CN_out_sig(2508);
VN_in_sig(3705)	<=	CN_out_sig(2509);
VN_in_sig(4213)	<=	CN_out_sig(2510);
VN_in_sig(4833)	<=	CN_out_sig(2511);
VN_in_sig(489)	<=	CN_out_sig(2512);
VN_in_sig(1081)	<=	CN_out_sig(2513);
VN_in_sig(1729)	<=	CN_out_sig(2514);
VN_in_sig(2193)	<=	CN_out_sig(2515);
VN_in_sig(2777)	<=	CN_out_sig(2516);
VN_in_sig(3709)	<=	CN_out_sig(2517);
VN_in_sig(4217)	<=	CN_out_sig(2518);
VN_in_sig(4837)	<=	CN_out_sig(2519);
VN_in_sig(493)	<=	CN_out_sig(2520);
VN_in_sig(1085)	<=	CN_out_sig(2521);
VN_in_sig(1733)	<=	CN_out_sig(2522);
VN_in_sig(2197)	<=	CN_out_sig(2523);
VN_in_sig(2781)	<=	CN_out_sig(2524);
VN_in_sig(3713)	<=	CN_out_sig(2525);
VN_in_sig(4221)	<=	CN_out_sig(2526);
VN_in_sig(4841)	<=	CN_out_sig(2527);
VN_in_sig(497)	<=	CN_out_sig(2528);
VN_in_sig(1089)	<=	CN_out_sig(2529);
VN_in_sig(1737)	<=	CN_out_sig(2530);
VN_in_sig(2201)	<=	CN_out_sig(2531);
VN_in_sig(2785)	<=	CN_out_sig(2532);
VN_in_sig(3717)	<=	CN_out_sig(2533);
VN_in_sig(4225)	<=	CN_out_sig(2534);
VN_in_sig(4845)	<=	CN_out_sig(2535);
VN_in_sig(501)	<=	CN_out_sig(2536);
VN_in_sig(1093)	<=	CN_out_sig(2537);
VN_in_sig(1741)	<=	CN_out_sig(2538);
VN_in_sig(2205)	<=	CN_out_sig(2539);
VN_in_sig(2789)	<=	CN_out_sig(2540);
VN_in_sig(3721)	<=	CN_out_sig(2541);
VN_in_sig(4229)	<=	CN_out_sig(2542);
VN_in_sig(4849)	<=	CN_out_sig(2543);
VN_in_sig(505)	<=	CN_out_sig(2544);
VN_in_sig(1097)	<=	CN_out_sig(2545);
VN_in_sig(1745)	<=	CN_out_sig(2546);
VN_in_sig(2209)	<=	CN_out_sig(2547);
VN_in_sig(2793)	<=	CN_out_sig(2548);
VN_in_sig(3725)	<=	CN_out_sig(2549);
VN_in_sig(4233)	<=	CN_out_sig(2550);
VN_in_sig(4853)	<=	CN_out_sig(2551);
VN_in_sig(509)	<=	CN_out_sig(2552);
VN_in_sig(1101)	<=	CN_out_sig(2553);
VN_in_sig(1749)	<=	CN_out_sig(2554);
VN_in_sig(2213)	<=	CN_out_sig(2555);
VN_in_sig(2797)	<=	CN_out_sig(2556);
VN_in_sig(3729)	<=	CN_out_sig(2557);
VN_in_sig(4237)	<=	CN_out_sig(2558);
VN_in_sig(4857)	<=	CN_out_sig(2559);
VN_in_sig(513)	<=	CN_out_sig(2560);
VN_in_sig(1105)	<=	CN_out_sig(2561);
VN_in_sig(1753)	<=	CN_out_sig(2562);
VN_in_sig(2217)	<=	CN_out_sig(2563);
VN_in_sig(2801)	<=	CN_out_sig(2564);
VN_in_sig(3733)	<=	CN_out_sig(2565);
VN_in_sig(4241)	<=	CN_out_sig(2566);
VN_in_sig(4861)	<=	CN_out_sig(2567);
VN_in_sig(517)	<=	CN_out_sig(2568);
VN_in_sig(1109)	<=	CN_out_sig(2569);
VN_in_sig(1757)	<=	CN_out_sig(2570);
VN_in_sig(2221)	<=	CN_out_sig(2571);
VN_in_sig(2805)	<=	CN_out_sig(2572);
VN_in_sig(3737)	<=	CN_out_sig(2573);
VN_in_sig(4245)	<=	CN_out_sig(2574);
VN_in_sig(4865)	<=	CN_out_sig(2575);
VN_in_sig(521)	<=	CN_out_sig(2576);
VN_in_sig(1113)	<=	CN_out_sig(2577);
VN_in_sig(1761)	<=	CN_out_sig(2578);
VN_in_sig(2225)	<=	CN_out_sig(2579);
VN_in_sig(2593)	<=	CN_out_sig(2580);
VN_in_sig(3741)	<=	CN_out_sig(2581);
VN_in_sig(4249)	<=	CN_out_sig(2582);
VN_in_sig(4869)	<=	CN_out_sig(2583);
VN_in_sig(525)	<=	CN_out_sig(2584);
VN_in_sig(1117)	<=	CN_out_sig(2585);
VN_in_sig(1765)	<=	CN_out_sig(2586);
VN_in_sig(2229)	<=	CN_out_sig(2587);
VN_in_sig(2597)	<=	CN_out_sig(2588);
VN_in_sig(3745)	<=	CN_out_sig(2589);
VN_in_sig(4253)	<=	CN_out_sig(2590);
VN_in_sig(4873)	<=	CN_out_sig(2591);
VN_in_sig(594)	<=	CN_out_sig(2592);
VN_in_sig(1222)	<=	CN_out_sig(2593);
VN_in_sig(1854)	<=	CN_out_sig(2594);
VN_in_sig(2022)	<=	CN_out_sig(2595);
VN_in_sig(2606)	<=	CN_out_sig(2596);
VN_in_sig(3410)	<=	CN_out_sig(2597);
VN_in_sig(4274)	<=	CN_out_sig(2598);
VN_in_sig(4910)	<=	CN_out_sig(2599);
VN_in_sig(598)	<=	CN_out_sig(2600);
VN_in_sig(1226)	<=	CN_out_sig(2601);
VN_in_sig(1858)	<=	CN_out_sig(2602);
VN_in_sig(2026)	<=	CN_out_sig(2603);
VN_in_sig(2610)	<=	CN_out_sig(2604);
VN_in_sig(3414)	<=	CN_out_sig(2605);
VN_in_sig(4278)	<=	CN_out_sig(2606);
VN_in_sig(4914)	<=	CN_out_sig(2607);
VN_in_sig(602)	<=	CN_out_sig(2608);
VN_in_sig(1230)	<=	CN_out_sig(2609);
VN_in_sig(1862)	<=	CN_out_sig(2610);
VN_in_sig(2030)	<=	CN_out_sig(2611);
VN_in_sig(2614)	<=	CN_out_sig(2612);
VN_in_sig(3418)	<=	CN_out_sig(2613);
VN_in_sig(4282)	<=	CN_out_sig(2614);
VN_in_sig(4918)	<=	CN_out_sig(2615);
VN_in_sig(606)	<=	CN_out_sig(2616);
VN_in_sig(1234)	<=	CN_out_sig(2617);
VN_in_sig(1866)	<=	CN_out_sig(2618);
VN_in_sig(2034)	<=	CN_out_sig(2619);
VN_in_sig(2618)	<=	CN_out_sig(2620);
VN_in_sig(3422)	<=	CN_out_sig(2621);
VN_in_sig(4286)	<=	CN_out_sig(2622);
VN_in_sig(4922)	<=	CN_out_sig(2623);
VN_in_sig(610)	<=	CN_out_sig(2624);
VN_in_sig(1238)	<=	CN_out_sig(2625);
VN_in_sig(1870)	<=	CN_out_sig(2626);
VN_in_sig(2038)	<=	CN_out_sig(2627);
VN_in_sig(2622)	<=	CN_out_sig(2628);
VN_in_sig(3426)	<=	CN_out_sig(2629);
VN_in_sig(4290)	<=	CN_out_sig(2630);
VN_in_sig(4926)	<=	CN_out_sig(2631);
VN_in_sig(614)	<=	CN_out_sig(2632);
VN_in_sig(1242)	<=	CN_out_sig(2633);
VN_in_sig(1874)	<=	CN_out_sig(2634);
VN_in_sig(2042)	<=	CN_out_sig(2635);
VN_in_sig(2626)	<=	CN_out_sig(2636);
VN_in_sig(3430)	<=	CN_out_sig(2637);
VN_in_sig(4294)	<=	CN_out_sig(2638);
VN_in_sig(4930)	<=	CN_out_sig(2639);
VN_in_sig(618)	<=	CN_out_sig(2640);
VN_in_sig(1246)	<=	CN_out_sig(2641);
VN_in_sig(1878)	<=	CN_out_sig(2642);
VN_in_sig(2046)	<=	CN_out_sig(2643);
VN_in_sig(2630)	<=	CN_out_sig(2644);
VN_in_sig(3434)	<=	CN_out_sig(2645);
VN_in_sig(4298)	<=	CN_out_sig(2646);
VN_in_sig(4934)	<=	CN_out_sig(2647);
VN_in_sig(622)	<=	CN_out_sig(2648);
VN_in_sig(1250)	<=	CN_out_sig(2649);
VN_in_sig(1882)	<=	CN_out_sig(2650);
VN_in_sig(2050)	<=	CN_out_sig(2651);
VN_in_sig(2634)	<=	CN_out_sig(2652);
VN_in_sig(3438)	<=	CN_out_sig(2653);
VN_in_sig(4302)	<=	CN_out_sig(2654);
VN_in_sig(4938)	<=	CN_out_sig(2655);
VN_in_sig(626)	<=	CN_out_sig(2656);
VN_in_sig(1254)	<=	CN_out_sig(2657);
VN_in_sig(1886)	<=	CN_out_sig(2658);
VN_in_sig(2054)	<=	CN_out_sig(2659);
VN_in_sig(2638)	<=	CN_out_sig(2660);
VN_in_sig(3442)	<=	CN_out_sig(2661);
VN_in_sig(4306)	<=	CN_out_sig(2662);
VN_in_sig(4942)	<=	CN_out_sig(2663);
VN_in_sig(630)	<=	CN_out_sig(2664);
VN_in_sig(1258)	<=	CN_out_sig(2665);
VN_in_sig(1890)	<=	CN_out_sig(2666);
VN_in_sig(2058)	<=	CN_out_sig(2667);
VN_in_sig(2642)	<=	CN_out_sig(2668);
VN_in_sig(3446)	<=	CN_out_sig(2669);
VN_in_sig(4310)	<=	CN_out_sig(2670);
VN_in_sig(4946)	<=	CN_out_sig(2671);
VN_in_sig(634)	<=	CN_out_sig(2672);
VN_in_sig(1262)	<=	CN_out_sig(2673);
VN_in_sig(1894)	<=	CN_out_sig(2674);
VN_in_sig(2062)	<=	CN_out_sig(2675);
VN_in_sig(2646)	<=	CN_out_sig(2676);
VN_in_sig(3450)	<=	CN_out_sig(2677);
VN_in_sig(4314)	<=	CN_out_sig(2678);
VN_in_sig(4950)	<=	CN_out_sig(2679);
VN_in_sig(638)	<=	CN_out_sig(2680);
VN_in_sig(1266)	<=	CN_out_sig(2681);
VN_in_sig(1898)	<=	CN_out_sig(2682);
VN_in_sig(2066)	<=	CN_out_sig(2683);
VN_in_sig(2650)	<=	CN_out_sig(2684);
VN_in_sig(3454)	<=	CN_out_sig(2685);
VN_in_sig(4318)	<=	CN_out_sig(2686);
VN_in_sig(4954)	<=	CN_out_sig(2687);
VN_in_sig(642)	<=	CN_out_sig(2688);
VN_in_sig(1270)	<=	CN_out_sig(2689);
VN_in_sig(1902)	<=	CN_out_sig(2690);
VN_in_sig(2070)	<=	CN_out_sig(2691);
VN_in_sig(2654)	<=	CN_out_sig(2692);
VN_in_sig(3242)	<=	CN_out_sig(2693);
VN_in_sig(4106)	<=	CN_out_sig(2694);
VN_in_sig(4958)	<=	CN_out_sig(2695);
VN_in_sig(646)	<=	CN_out_sig(2696);
VN_in_sig(1274)	<=	CN_out_sig(2697);
VN_in_sig(1906)	<=	CN_out_sig(2698);
VN_in_sig(2074)	<=	CN_out_sig(2699);
VN_in_sig(2658)	<=	CN_out_sig(2700);
VN_in_sig(3246)	<=	CN_out_sig(2701);
VN_in_sig(4110)	<=	CN_out_sig(2702);
VN_in_sig(4962)	<=	CN_out_sig(2703);
VN_in_sig(434)	<=	CN_out_sig(2704);
VN_in_sig(1278)	<=	CN_out_sig(2705);
VN_in_sig(1910)	<=	CN_out_sig(2706);
VN_in_sig(2078)	<=	CN_out_sig(2707);
VN_in_sig(2662)	<=	CN_out_sig(2708);
VN_in_sig(3250)	<=	CN_out_sig(2709);
VN_in_sig(4114)	<=	CN_out_sig(2710);
VN_in_sig(4966)	<=	CN_out_sig(2711);
VN_in_sig(438)	<=	CN_out_sig(2712);
VN_in_sig(1282)	<=	CN_out_sig(2713);
VN_in_sig(1914)	<=	CN_out_sig(2714);
VN_in_sig(2082)	<=	CN_out_sig(2715);
VN_in_sig(2666)	<=	CN_out_sig(2716);
VN_in_sig(3254)	<=	CN_out_sig(2717);
VN_in_sig(4118)	<=	CN_out_sig(2718);
VN_in_sig(4754)	<=	CN_out_sig(2719);
VN_in_sig(442)	<=	CN_out_sig(2720);
VN_in_sig(1286)	<=	CN_out_sig(2721);
VN_in_sig(1918)	<=	CN_out_sig(2722);
VN_in_sig(2086)	<=	CN_out_sig(2723);
VN_in_sig(2670)	<=	CN_out_sig(2724);
VN_in_sig(3258)	<=	CN_out_sig(2725);
VN_in_sig(4122)	<=	CN_out_sig(2726);
VN_in_sig(4758)	<=	CN_out_sig(2727);
VN_in_sig(446)	<=	CN_out_sig(2728);
VN_in_sig(1290)	<=	CN_out_sig(2729);
VN_in_sig(1922)	<=	CN_out_sig(2730);
VN_in_sig(2090)	<=	CN_out_sig(2731);
VN_in_sig(2674)	<=	CN_out_sig(2732);
VN_in_sig(3262)	<=	CN_out_sig(2733);
VN_in_sig(4126)	<=	CN_out_sig(2734);
VN_in_sig(4762)	<=	CN_out_sig(2735);
VN_in_sig(450)	<=	CN_out_sig(2736);
VN_in_sig(1294)	<=	CN_out_sig(2737);
VN_in_sig(1926)	<=	CN_out_sig(2738);
VN_in_sig(2094)	<=	CN_out_sig(2739);
VN_in_sig(2678)	<=	CN_out_sig(2740);
VN_in_sig(3266)	<=	CN_out_sig(2741);
VN_in_sig(4130)	<=	CN_out_sig(2742);
VN_in_sig(4766)	<=	CN_out_sig(2743);
VN_in_sig(454)	<=	CN_out_sig(2744);
VN_in_sig(1082)	<=	CN_out_sig(2745);
VN_in_sig(1930)	<=	CN_out_sig(2746);
VN_in_sig(2098)	<=	CN_out_sig(2747);
VN_in_sig(2682)	<=	CN_out_sig(2748);
VN_in_sig(3270)	<=	CN_out_sig(2749);
VN_in_sig(4134)	<=	CN_out_sig(2750);
VN_in_sig(4770)	<=	CN_out_sig(2751);
VN_in_sig(458)	<=	CN_out_sig(2752);
VN_in_sig(1086)	<=	CN_out_sig(2753);
VN_in_sig(1934)	<=	CN_out_sig(2754);
VN_in_sig(2102)	<=	CN_out_sig(2755);
VN_in_sig(2686)	<=	CN_out_sig(2756);
VN_in_sig(3274)	<=	CN_out_sig(2757);
VN_in_sig(4138)	<=	CN_out_sig(2758);
VN_in_sig(4774)	<=	CN_out_sig(2759);
VN_in_sig(462)	<=	CN_out_sig(2760);
VN_in_sig(1090)	<=	CN_out_sig(2761);
VN_in_sig(1938)	<=	CN_out_sig(2762);
VN_in_sig(2106)	<=	CN_out_sig(2763);
VN_in_sig(2690)	<=	CN_out_sig(2764);
VN_in_sig(3278)	<=	CN_out_sig(2765);
VN_in_sig(4142)	<=	CN_out_sig(2766);
VN_in_sig(4778)	<=	CN_out_sig(2767);
VN_in_sig(466)	<=	CN_out_sig(2768);
VN_in_sig(1094)	<=	CN_out_sig(2769);
VN_in_sig(1942)	<=	CN_out_sig(2770);
VN_in_sig(2110)	<=	CN_out_sig(2771);
VN_in_sig(2694)	<=	CN_out_sig(2772);
VN_in_sig(3282)	<=	CN_out_sig(2773);
VN_in_sig(4146)	<=	CN_out_sig(2774);
VN_in_sig(4782)	<=	CN_out_sig(2775);
VN_in_sig(470)	<=	CN_out_sig(2776);
VN_in_sig(1098)	<=	CN_out_sig(2777);
VN_in_sig(1730)	<=	CN_out_sig(2778);
VN_in_sig(2114)	<=	CN_out_sig(2779);
VN_in_sig(2698)	<=	CN_out_sig(2780);
VN_in_sig(3286)	<=	CN_out_sig(2781);
VN_in_sig(4150)	<=	CN_out_sig(2782);
VN_in_sig(4786)	<=	CN_out_sig(2783);
VN_in_sig(474)	<=	CN_out_sig(2784);
VN_in_sig(1102)	<=	CN_out_sig(2785);
VN_in_sig(1734)	<=	CN_out_sig(2786);
VN_in_sig(2118)	<=	CN_out_sig(2787);
VN_in_sig(2702)	<=	CN_out_sig(2788);
VN_in_sig(3290)	<=	CN_out_sig(2789);
VN_in_sig(4154)	<=	CN_out_sig(2790);
VN_in_sig(4790)	<=	CN_out_sig(2791);
VN_in_sig(478)	<=	CN_out_sig(2792);
VN_in_sig(1106)	<=	CN_out_sig(2793);
VN_in_sig(1738)	<=	CN_out_sig(2794);
VN_in_sig(2122)	<=	CN_out_sig(2795);
VN_in_sig(2706)	<=	CN_out_sig(2796);
VN_in_sig(3294)	<=	CN_out_sig(2797);
VN_in_sig(4158)	<=	CN_out_sig(2798);
VN_in_sig(4794)	<=	CN_out_sig(2799);
VN_in_sig(482)	<=	CN_out_sig(2800);
VN_in_sig(1110)	<=	CN_out_sig(2801);
VN_in_sig(1742)	<=	CN_out_sig(2802);
VN_in_sig(2126)	<=	CN_out_sig(2803);
VN_in_sig(2710)	<=	CN_out_sig(2804);
VN_in_sig(3298)	<=	CN_out_sig(2805);
VN_in_sig(4162)	<=	CN_out_sig(2806);
VN_in_sig(4798)	<=	CN_out_sig(2807);
VN_in_sig(486)	<=	CN_out_sig(2808);
VN_in_sig(1114)	<=	CN_out_sig(2809);
VN_in_sig(1746)	<=	CN_out_sig(2810);
VN_in_sig(2130)	<=	CN_out_sig(2811);
VN_in_sig(2714)	<=	CN_out_sig(2812);
VN_in_sig(3302)	<=	CN_out_sig(2813);
VN_in_sig(4166)	<=	CN_out_sig(2814);
VN_in_sig(4802)	<=	CN_out_sig(2815);
VN_in_sig(490)	<=	CN_out_sig(2816);
VN_in_sig(1118)	<=	CN_out_sig(2817);
VN_in_sig(1750)	<=	CN_out_sig(2818);
VN_in_sig(2134)	<=	CN_out_sig(2819);
VN_in_sig(2718)	<=	CN_out_sig(2820);
VN_in_sig(3306)	<=	CN_out_sig(2821);
VN_in_sig(4170)	<=	CN_out_sig(2822);
VN_in_sig(4806)	<=	CN_out_sig(2823);
VN_in_sig(494)	<=	CN_out_sig(2824);
VN_in_sig(1122)	<=	CN_out_sig(2825);
VN_in_sig(1754)	<=	CN_out_sig(2826);
VN_in_sig(2138)	<=	CN_out_sig(2827);
VN_in_sig(2722)	<=	CN_out_sig(2828);
VN_in_sig(3310)	<=	CN_out_sig(2829);
VN_in_sig(4174)	<=	CN_out_sig(2830);
VN_in_sig(4810)	<=	CN_out_sig(2831);
VN_in_sig(498)	<=	CN_out_sig(2832);
VN_in_sig(1126)	<=	CN_out_sig(2833);
VN_in_sig(1758)	<=	CN_out_sig(2834);
VN_in_sig(2142)	<=	CN_out_sig(2835);
VN_in_sig(2726)	<=	CN_out_sig(2836);
VN_in_sig(3314)	<=	CN_out_sig(2837);
VN_in_sig(4178)	<=	CN_out_sig(2838);
VN_in_sig(4814)	<=	CN_out_sig(2839);
VN_in_sig(502)	<=	CN_out_sig(2840);
VN_in_sig(1130)	<=	CN_out_sig(2841);
VN_in_sig(1762)	<=	CN_out_sig(2842);
VN_in_sig(2146)	<=	CN_out_sig(2843);
VN_in_sig(2730)	<=	CN_out_sig(2844);
VN_in_sig(3318)	<=	CN_out_sig(2845);
VN_in_sig(4182)	<=	CN_out_sig(2846);
VN_in_sig(4818)	<=	CN_out_sig(2847);
VN_in_sig(506)	<=	CN_out_sig(2848);
VN_in_sig(1134)	<=	CN_out_sig(2849);
VN_in_sig(1766)	<=	CN_out_sig(2850);
VN_in_sig(2150)	<=	CN_out_sig(2851);
VN_in_sig(2734)	<=	CN_out_sig(2852);
VN_in_sig(3322)	<=	CN_out_sig(2853);
VN_in_sig(4186)	<=	CN_out_sig(2854);
VN_in_sig(4822)	<=	CN_out_sig(2855);
VN_in_sig(510)	<=	CN_out_sig(2856);
VN_in_sig(1138)	<=	CN_out_sig(2857);
VN_in_sig(1770)	<=	CN_out_sig(2858);
VN_in_sig(2154)	<=	CN_out_sig(2859);
VN_in_sig(2738)	<=	CN_out_sig(2860);
VN_in_sig(3326)	<=	CN_out_sig(2861);
VN_in_sig(4190)	<=	CN_out_sig(2862);
VN_in_sig(4826)	<=	CN_out_sig(2863);
VN_in_sig(514)	<=	CN_out_sig(2864);
VN_in_sig(1142)	<=	CN_out_sig(2865);
VN_in_sig(1774)	<=	CN_out_sig(2866);
VN_in_sig(2158)	<=	CN_out_sig(2867);
VN_in_sig(2742)	<=	CN_out_sig(2868);
VN_in_sig(3330)	<=	CN_out_sig(2869);
VN_in_sig(4194)	<=	CN_out_sig(2870);
VN_in_sig(4830)	<=	CN_out_sig(2871);
VN_in_sig(518)	<=	CN_out_sig(2872);
VN_in_sig(1146)	<=	CN_out_sig(2873);
VN_in_sig(1778)	<=	CN_out_sig(2874);
VN_in_sig(1946)	<=	CN_out_sig(2875);
VN_in_sig(2746)	<=	CN_out_sig(2876);
VN_in_sig(3334)	<=	CN_out_sig(2877);
VN_in_sig(4198)	<=	CN_out_sig(2878);
VN_in_sig(4834)	<=	CN_out_sig(2879);
VN_in_sig(522)	<=	CN_out_sig(2880);
VN_in_sig(1150)	<=	CN_out_sig(2881);
VN_in_sig(1782)	<=	CN_out_sig(2882);
VN_in_sig(1950)	<=	CN_out_sig(2883);
VN_in_sig(2750)	<=	CN_out_sig(2884);
VN_in_sig(3338)	<=	CN_out_sig(2885);
VN_in_sig(4202)	<=	CN_out_sig(2886);
VN_in_sig(4838)	<=	CN_out_sig(2887);
VN_in_sig(526)	<=	CN_out_sig(2888);
VN_in_sig(1154)	<=	CN_out_sig(2889);
VN_in_sig(1786)	<=	CN_out_sig(2890);
VN_in_sig(1954)	<=	CN_out_sig(2891);
VN_in_sig(2754)	<=	CN_out_sig(2892);
VN_in_sig(3342)	<=	CN_out_sig(2893);
VN_in_sig(4206)	<=	CN_out_sig(2894);
VN_in_sig(4842)	<=	CN_out_sig(2895);
VN_in_sig(530)	<=	CN_out_sig(2896);
VN_in_sig(1158)	<=	CN_out_sig(2897);
VN_in_sig(1790)	<=	CN_out_sig(2898);
VN_in_sig(1958)	<=	CN_out_sig(2899);
VN_in_sig(2758)	<=	CN_out_sig(2900);
VN_in_sig(3346)	<=	CN_out_sig(2901);
VN_in_sig(4210)	<=	CN_out_sig(2902);
VN_in_sig(4846)	<=	CN_out_sig(2903);
VN_in_sig(534)	<=	CN_out_sig(2904);
VN_in_sig(1162)	<=	CN_out_sig(2905);
VN_in_sig(1794)	<=	CN_out_sig(2906);
VN_in_sig(1962)	<=	CN_out_sig(2907);
VN_in_sig(2762)	<=	CN_out_sig(2908);
VN_in_sig(3350)	<=	CN_out_sig(2909);
VN_in_sig(4214)	<=	CN_out_sig(2910);
VN_in_sig(4850)	<=	CN_out_sig(2911);
VN_in_sig(538)	<=	CN_out_sig(2912);
VN_in_sig(1166)	<=	CN_out_sig(2913);
VN_in_sig(1798)	<=	CN_out_sig(2914);
VN_in_sig(1966)	<=	CN_out_sig(2915);
VN_in_sig(2766)	<=	CN_out_sig(2916);
VN_in_sig(3354)	<=	CN_out_sig(2917);
VN_in_sig(4218)	<=	CN_out_sig(2918);
VN_in_sig(4854)	<=	CN_out_sig(2919);
VN_in_sig(542)	<=	CN_out_sig(2920);
VN_in_sig(1170)	<=	CN_out_sig(2921);
VN_in_sig(1802)	<=	CN_out_sig(2922);
VN_in_sig(1970)	<=	CN_out_sig(2923);
VN_in_sig(2770)	<=	CN_out_sig(2924);
VN_in_sig(3358)	<=	CN_out_sig(2925);
VN_in_sig(4222)	<=	CN_out_sig(2926);
VN_in_sig(4858)	<=	CN_out_sig(2927);
VN_in_sig(546)	<=	CN_out_sig(2928);
VN_in_sig(1174)	<=	CN_out_sig(2929);
VN_in_sig(1806)	<=	CN_out_sig(2930);
VN_in_sig(1974)	<=	CN_out_sig(2931);
VN_in_sig(2774)	<=	CN_out_sig(2932);
VN_in_sig(3362)	<=	CN_out_sig(2933);
VN_in_sig(4226)	<=	CN_out_sig(2934);
VN_in_sig(4862)	<=	CN_out_sig(2935);
VN_in_sig(550)	<=	CN_out_sig(2936);
VN_in_sig(1178)	<=	CN_out_sig(2937);
VN_in_sig(1810)	<=	CN_out_sig(2938);
VN_in_sig(1978)	<=	CN_out_sig(2939);
VN_in_sig(2778)	<=	CN_out_sig(2940);
VN_in_sig(3366)	<=	CN_out_sig(2941);
VN_in_sig(4230)	<=	CN_out_sig(2942);
VN_in_sig(4866)	<=	CN_out_sig(2943);
VN_in_sig(554)	<=	CN_out_sig(2944);
VN_in_sig(1182)	<=	CN_out_sig(2945);
VN_in_sig(1814)	<=	CN_out_sig(2946);
VN_in_sig(1982)	<=	CN_out_sig(2947);
VN_in_sig(2782)	<=	CN_out_sig(2948);
VN_in_sig(3370)	<=	CN_out_sig(2949);
VN_in_sig(4234)	<=	CN_out_sig(2950);
VN_in_sig(4870)	<=	CN_out_sig(2951);
VN_in_sig(558)	<=	CN_out_sig(2952);
VN_in_sig(1186)	<=	CN_out_sig(2953);
VN_in_sig(1818)	<=	CN_out_sig(2954);
VN_in_sig(1986)	<=	CN_out_sig(2955);
VN_in_sig(2786)	<=	CN_out_sig(2956);
VN_in_sig(3374)	<=	CN_out_sig(2957);
VN_in_sig(4238)	<=	CN_out_sig(2958);
VN_in_sig(4874)	<=	CN_out_sig(2959);
VN_in_sig(562)	<=	CN_out_sig(2960);
VN_in_sig(1190)	<=	CN_out_sig(2961);
VN_in_sig(1822)	<=	CN_out_sig(2962);
VN_in_sig(1990)	<=	CN_out_sig(2963);
VN_in_sig(2790)	<=	CN_out_sig(2964);
VN_in_sig(3378)	<=	CN_out_sig(2965);
VN_in_sig(4242)	<=	CN_out_sig(2966);
VN_in_sig(4878)	<=	CN_out_sig(2967);
VN_in_sig(566)	<=	CN_out_sig(2968);
VN_in_sig(1194)	<=	CN_out_sig(2969);
VN_in_sig(1826)	<=	CN_out_sig(2970);
VN_in_sig(1994)	<=	CN_out_sig(2971);
VN_in_sig(2794)	<=	CN_out_sig(2972);
VN_in_sig(3382)	<=	CN_out_sig(2973);
VN_in_sig(4246)	<=	CN_out_sig(2974);
VN_in_sig(4882)	<=	CN_out_sig(2975);
VN_in_sig(570)	<=	CN_out_sig(2976);
VN_in_sig(1198)	<=	CN_out_sig(2977);
VN_in_sig(1830)	<=	CN_out_sig(2978);
VN_in_sig(1998)	<=	CN_out_sig(2979);
VN_in_sig(2798)	<=	CN_out_sig(2980);
VN_in_sig(3386)	<=	CN_out_sig(2981);
VN_in_sig(4250)	<=	CN_out_sig(2982);
VN_in_sig(4886)	<=	CN_out_sig(2983);
VN_in_sig(574)	<=	CN_out_sig(2984);
VN_in_sig(1202)	<=	CN_out_sig(2985);
VN_in_sig(1834)	<=	CN_out_sig(2986);
VN_in_sig(2002)	<=	CN_out_sig(2987);
VN_in_sig(2802)	<=	CN_out_sig(2988);
VN_in_sig(3390)	<=	CN_out_sig(2989);
VN_in_sig(4254)	<=	CN_out_sig(2990);
VN_in_sig(4890)	<=	CN_out_sig(2991);
VN_in_sig(578)	<=	CN_out_sig(2992);
VN_in_sig(1206)	<=	CN_out_sig(2993);
VN_in_sig(1838)	<=	CN_out_sig(2994);
VN_in_sig(2006)	<=	CN_out_sig(2995);
VN_in_sig(2806)	<=	CN_out_sig(2996);
VN_in_sig(3394)	<=	CN_out_sig(2997);
VN_in_sig(4258)	<=	CN_out_sig(2998);
VN_in_sig(4894)	<=	CN_out_sig(2999);
VN_in_sig(582)	<=	CN_out_sig(3000);
VN_in_sig(1210)	<=	CN_out_sig(3001);
VN_in_sig(1842)	<=	CN_out_sig(3002);
VN_in_sig(2010)	<=	CN_out_sig(3003);
VN_in_sig(2594)	<=	CN_out_sig(3004);
VN_in_sig(3398)	<=	CN_out_sig(3005);
VN_in_sig(4262)	<=	CN_out_sig(3006);
VN_in_sig(4898)	<=	CN_out_sig(3007);
VN_in_sig(586)	<=	CN_out_sig(3008);
VN_in_sig(1214)	<=	CN_out_sig(3009);
VN_in_sig(1846)	<=	CN_out_sig(3010);
VN_in_sig(2014)	<=	CN_out_sig(3011);
VN_in_sig(2598)	<=	CN_out_sig(3012);
VN_in_sig(3402)	<=	CN_out_sig(3013);
VN_in_sig(4266)	<=	CN_out_sig(3014);
VN_in_sig(4902)	<=	CN_out_sig(3015);
VN_in_sig(590)	<=	CN_out_sig(3016);
VN_in_sig(1218)	<=	CN_out_sig(3017);
VN_in_sig(1850)	<=	CN_out_sig(3018);
VN_in_sig(2018)	<=	CN_out_sig(3019);
VN_in_sig(2602)	<=	CN_out_sig(3020);
VN_in_sig(3406)	<=	CN_out_sig(3021);
VN_in_sig(4270)	<=	CN_out_sig(3022);
VN_in_sig(4906)	<=	CN_out_sig(3023);
VN_in_sig(334)	<=	CN_out_sig(3024);
VN_in_sig(650)	<=	CN_out_sig(3025);
VN_in_sig(1630)	<=	CN_out_sig(3026);
VN_in_sig(2182)	<=	CN_out_sig(3027);
VN_in_sig(3214)	<=	CN_out_sig(3028);
VN_in_sig(3786)	<=	CN_out_sig(3029);
VN_in_sig(4434)	<=	CN_out_sig(3030);
VN_in_sig(4702)	<=	CN_out_sig(3031);
VN_in_sig(338)	<=	CN_out_sig(3032);
VN_in_sig(654)	<=	CN_out_sig(3033);
VN_in_sig(1634)	<=	CN_out_sig(3034);
VN_in_sig(2186)	<=	CN_out_sig(3035);
VN_in_sig(3218)	<=	CN_out_sig(3036);
VN_in_sig(3790)	<=	CN_out_sig(3037);
VN_in_sig(4438)	<=	CN_out_sig(3038);
VN_in_sig(4706)	<=	CN_out_sig(3039);
VN_in_sig(342)	<=	CN_out_sig(3040);
VN_in_sig(658)	<=	CN_out_sig(3041);
VN_in_sig(1638)	<=	CN_out_sig(3042);
VN_in_sig(2190)	<=	CN_out_sig(3043);
VN_in_sig(3222)	<=	CN_out_sig(3044);
VN_in_sig(3794)	<=	CN_out_sig(3045);
VN_in_sig(4442)	<=	CN_out_sig(3046);
VN_in_sig(4710)	<=	CN_out_sig(3047);
VN_in_sig(346)	<=	CN_out_sig(3048);
VN_in_sig(662)	<=	CN_out_sig(3049);
VN_in_sig(1642)	<=	CN_out_sig(3050);
VN_in_sig(2194)	<=	CN_out_sig(3051);
VN_in_sig(3226)	<=	CN_out_sig(3052);
VN_in_sig(3798)	<=	CN_out_sig(3053);
VN_in_sig(4446)	<=	CN_out_sig(3054);
VN_in_sig(4714)	<=	CN_out_sig(3055);
VN_in_sig(350)	<=	CN_out_sig(3056);
VN_in_sig(666)	<=	CN_out_sig(3057);
VN_in_sig(1646)	<=	CN_out_sig(3058);
VN_in_sig(2198)	<=	CN_out_sig(3059);
VN_in_sig(3230)	<=	CN_out_sig(3060);
VN_in_sig(3802)	<=	CN_out_sig(3061);
VN_in_sig(4450)	<=	CN_out_sig(3062);
VN_in_sig(4718)	<=	CN_out_sig(3063);
VN_in_sig(354)	<=	CN_out_sig(3064);
VN_in_sig(670)	<=	CN_out_sig(3065);
VN_in_sig(1650)	<=	CN_out_sig(3066);
VN_in_sig(2202)	<=	CN_out_sig(3067);
VN_in_sig(3234)	<=	CN_out_sig(3068);
VN_in_sig(3806)	<=	CN_out_sig(3069);
VN_in_sig(4454)	<=	CN_out_sig(3070);
VN_in_sig(4722)	<=	CN_out_sig(3071);
VN_in_sig(358)	<=	CN_out_sig(3072);
VN_in_sig(674)	<=	CN_out_sig(3073);
VN_in_sig(1654)	<=	CN_out_sig(3074);
VN_in_sig(2206)	<=	CN_out_sig(3075);
VN_in_sig(3238)	<=	CN_out_sig(3076);
VN_in_sig(3810)	<=	CN_out_sig(3077);
VN_in_sig(4458)	<=	CN_out_sig(3078);
VN_in_sig(4726)	<=	CN_out_sig(3079);
VN_in_sig(362)	<=	CN_out_sig(3080);
VN_in_sig(678)	<=	CN_out_sig(3081);
VN_in_sig(1658)	<=	CN_out_sig(3082);
VN_in_sig(2210)	<=	CN_out_sig(3083);
VN_in_sig(3026)	<=	CN_out_sig(3084);
VN_in_sig(3814)	<=	CN_out_sig(3085);
VN_in_sig(4462)	<=	CN_out_sig(3086);
VN_in_sig(4730)	<=	CN_out_sig(3087);
VN_in_sig(366)	<=	CN_out_sig(3088);
VN_in_sig(682)	<=	CN_out_sig(3089);
VN_in_sig(1662)	<=	CN_out_sig(3090);
VN_in_sig(2214)	<=	CN_out_sig(3091);
VN_in_sig(3030)	<=	CN_out_sig(3092);
VN_in_sig(3818)	<=	CN_out_sig(3093);
VN_in_sig(4466)	<=	CN_out_sig(3094);
VN_in_sig(4734)	<=	CN_out_sig(3095);
VN_in_sig(370)	<=	CN_out_sig(3096);
VN_in_sig(686)	<=	CN_out_sig(3097);
VN_in_sig(1666)	<=	CN_out_sig(3098);
VN_in_sig(2218)	<=	CN_out_sig(3099);
VN_in_sig(3034)	<=	CN_out_sig(3100);
VN_in_sig(3822)	<=	CN_out_sig(3101);
VN_in_sig(4470)	<=	CN_out_sig(3102);
VN_in_sig(4738)	<=	CN_out_sig(3103);
VN_in_sig(374)	<=	CN_out_sig(3104);
VN_in_sig(690)	<=	CN_out_sig(3105);
VN_in_sig(1670)	<=	CN_out_sig(3106);
VN_in_sig(2222)	<=	CN_out_sig(3107);
VN_in_sig(3038)	<=	CN_out_sig(3108);
VN_in_sig(3826)	<=	CN_out_sig(3109);
VN_in_sig(4474)	<=	CN_out_sig(3110);
VN_in_sig(4742)	<=	CN_out_sig(3111);
VN_in_sig(378)	<=	CN_out_sig(3112);
VN_in_sig(694)	<=	CN_out_sig(3113);
VN_in_sig(1674)	<=	CN_out_sig(3114);
VN_in_sig(2226)	<=	CN_out_sig(3115);
VN_in_sig(3042)	<=	CN_out_sig(3116);
VN_in_sig(3830)	<=	CN_out_sig(3117);
VN_in_sig(4478)	<=	CN_out_sig(3118);
VN_in_sig(4746)	<=	CN_out_sig(3119);
VN_in_sig(382)	<=	CN_out_sig(3120);
VN_in_sig(698)	<=	CN_out_sig(3121);
VN_in_sig(1678)	<=	CN_out_sig(3122);
VN_in_sig(2230)	<=	CN_out_sig(3123);
VN_in_sig(3046)	<=	CN_out_sig(3124);
VN_in_sig(3834)	<=	CN_out_sig(3125);
VN_in_sig(4482)	<=	CN_out_sig(3126);
VN_in_sig(4750)	<=	CN_out_sig(3127);
VN_in_sig(386)	<=	CN_out_sig(3128);
VN_in_sig(702)	<=	CN_out_sig(3129);
VN_in_sig(1682)	<=	CN_out_sig(3130);
VN_in_sig(2234)	<=	CN_out_sig(3131);
VN_in_sig(3050)	<=	CN_out_sig(3132);
VN_in_sig(3838)	<=	CN_out_sig(3133);
VN_in_sig(4486)	<=	CN_out_sig(3134);
VN_in_sig(4538)	<=	CN_out_sig(3135);
VN_in_sig(390)	<=	CN_out_sig(3136);
VN_in_sig(706)	<=	CN_out_sig(3137);
VN_in_sig(1686)	<=	CN_out_sig(3138);
VN_in_sig(2238)	<=	CN_out_sig(3139);
VN_in_sig(3054)	<=	CN_out_sig(3140);
VN_in_sig(3842)	<=	CN_out_sig(3141);
VN_in_sig(4490)	<=	CN_out_sig(3142);
VN_in_sig(4542)	<=	CN_out_sig(3143);
VN_in_sig(394)	<=	CN_out_sig(3144);
VN_in_sig(710)	<=	CN_out_sig(3145);
VN_in_sig(1690)	<=	CN_out_sig(3146);
VN_in_sig(2242)	<=	CN_out_sig(3147);
VN_in_sig(3058)	<=	CN_out_sig(3148);
VN_in_sig(3846)	<=	CN_out_sig(3149);
VN_in_sig(4494)	<=	CN_out_sig(3150);
VN_in_sig(4546)	<=	CN_out_sig(3151);
VN_in_sig(398)	<=	CN_out_sig(3152);
VN_in_sig(714)	<=	CN_out_sig(3153);
VN_in_sig(1694)	<=	CN_out_sig(3154);
VN_in_sig(2246)	<=	CN_out_sig(3155);
VN_in_sig(3062)	<=	CN_out_sig(3156);
VN_in_sig(3850)	<=	CN_out_sig(3157);
VN_in_sig(4498)	<=	CN_out_sig(3158);
VN_in_sig(4550)	<=	CN_out_sig(3159);
VN_in_sig(402)	<=	CN_out_sig(3160);
VN_in_sig(718)	<=	CN_out_sig(3161);
VN_in_sig(1698)	<=	CN_out_sig(3162);
VN_in_sig(2250)	<=	CN_out_sig(3163);
VN_in_sig(3066)	<=	CN_out_sig(3164);
VN_in_sig(3854)	<=	CN_out_sig(3165);
VN_in_sig(4502)	<=	CN_out_sig(3166);
VN_in_sig(4554)	<=	CN_out_sig(3167);
VN_in_sig(406)	<=	CN_out_sig(3168);
VN_in_sig(722)	<=	CN_out_sig(3169);
VN_in_sig(1702)	<=	CN_out_sig(3170);
VN_in_sig(2254)	<=	CN_out_sig(3171);
VN_in_sig(3070)	<=	CN_out_sig(3172);
VN_in_sig(3858)	<=	CN_out_sig(3173);
VN_in_sig(4506)	<=	CN_out_sig(3174);
VN_in_sig(4558)	<=	CN_out_sig(3175);
VN_in_sig(410)	<=	CN_out_sig(3176);
VN_in_sig(726)	<=	CN_out_sig(3177);
VN_in_sig(1706)	<=	CN_out_sig(3178);
VN_in_sig(2258)	<=	CN_out_sig(3179);
VN_in_sig(3074)	<=	CN_out_sig(3180);
VN_in_sig(3862)	<=	CN_out_sig(3181);
VN_in_sig(4510)	<=	CN_out_sig(3182);
VN_in_sig(4562)	<=	CN_out_sig(3183);
VN_in_sig(414)	<=	CN_out_sig(3184);
VN_in_sig(730)	<=	CN_out_sig(3185);
VN_in_sig(1710)	<=	CN_out_sig(3186);
VN_in_sig(2262)	<=	CN_out_sig(3187);
VN_in_sig(3078)	<=	CN_out_sig(3188);
VN_in_sig(3866)	<=	CN_out_sig(3189);
VN_in_sig(4514)	<=	CN_out_sig(3190);
VN_in_sig(4566)	<=	CN_out_sig(3191);
VN_in_sig(418)	<=	CN_out_sig(3192);
VN_in_sig(734)	<=	CN_out_sig(3193);
VN_in_sig(1714)	<=	CN_out_sig(3194);
VN_in_sig(2266)	<=	CN_out_sig(3195);
VN_in_sig(3082)	<=	CN_out_sig(3196);
VN_in_sig(3870)	<=	CN_out_sig(3197);
VN_in_sig(4518)	<=	CN_out_sig(3198);
VN_in_sig(4570)	<=	CN_out_sig(3199);
VN_in_sig(422)	<=	CN_out_sig(3200);
VN_in_sig(738)	<=	CN_out_sig(3201);
VN_in_sig(1718)	<=	CN_out_sig(3202);
VN_in_sig(2270)	<=	CN_out_sig(3203);
VN_in_sig(3086)	<=	CN_out_sig(3204);
VN_in_sig(3874)	<=	CN_out_sig(3205);
VN_in_sig(4522)	<=	CN_out_sig(3206);
VN_in_sig(4574)	<=	CN_out_sig(3207);
VN_in_sig(426)	<=	CN_out_sig(3208);
VN_in_sig(742)	<=	CN_out_sig(3209);
VN_in_sig(1722)	<=	CN_out_sig(3210);
VN_in_sig(2274)	<=	CN_out_sig(3211);
VN_in_sig(3090)	<=	CN_out_sig(3212);
VN_in_sig(3878)	<=	CN_out_sig(3213);
VN_in_sig(4526)	<=	CN_out_sig(3214);
VN_in_sig(4578)	<=	CN_out_sig(3215);
VN_in_sig(430)	<=	CN_out_sig(3216);
VN_in_sig(746)	<=	CN_out_sig(3217);
VN_in_sig(1726)	<=	CN_out_sig(3218);
VN_in_sig(2278)	<=	CN_out_sig(3219);
VN_in_sig(3094)	<=	CN_out_sig(3220);
VN_in_sig(3882)	<=	CN_out_sig(3221);
VN_in_sig(4530)	<=	CN_out_sig(3222);
VN_in_sig(4582)	<=	CN_out_sig(3223);
VN_in_sig(218)	<=	CN_out_sig(3224);
VN_in_sig(750)	<=	CN_out_sig(3225);
VN_in_sig(1514)	<=	CN_out_sig(3226);
VN_in_sig(2282)	<=	CN_out_sig(3227);
VN_in_sig(3098)	<=	CN_out_sig(3228);
VN_in_sig(3886)	<=	CN_out_sig(3229);
VN_in_sig(4534)	<=	CN_out_sig(3230);
VN_in_sig(4586)	<=	CN_out_sig(3231);
VN_in_sig(222)	<=	CN_out_sig(3232);
VN_in_sig(754)	<=	CN_out_sig(3233);
VN_in_sig(1518)	<=	CN_out_sig(3234);
VN_in_sig(2286)	<=	CN_out_sig(3235);
VN_in_sig(3102)	<=	CN_out_sig(3236);
VN_in_sig(3674)	<=	CN_out_sig(3237);
VN_in_sig(4322)	<=	CN_out_sig(3238);
VN_in_sig(4590)	<=	CN_out_sig(3239);
VN_in_sig(226)	<=	CN_out_sig(3240);
VN_in_sig(758)	<=	CN_out_sig(3241);
VN_in_sig(1522)	<=	CN_out_sig(3242);
VN_in_sig(2290)	<=	CN_out_sig(3243);
VN_in_sig(3106)	<=	CN_out_sig(3244);
VN_in_sig(3678)	<=	CN_out_sig(3245);
VN_in_sig(4326)	<=	CN_out_sig(3246);
VN_in_sig(4594)	<=	CN_out_sig(3247);
VN_in_sig(230)	<=	CN_out_sig(3248);
VN_in_sig(762)	<=	CN_out_sig(3249);
VN_in_sig(1526)	<=	CN_out_sig(3250);
VN_in_sig(2294)	<=	CN_out_sig(3251);
VN_in_sig(3110)	<=	CN_out_sig(3252);
VN_in_sig(3682)	<=	CN_out_sig(3253);
VN_in_sig(4330)	<=	CN_out_sig(3254);
VN_in_sig(4598)	<=	CN_out_sig(3255);
VN_in_sig(234)	<=	CN_out_sig(3256);
VN_in_sig(766)	<=	CN_out_sig(3257);
VN_in_sig(1530)	<=	CN_out_sig(3258);
VN_in_sig(2298)	<=	CN_out_sig(3259);
VN_in_sig(3114)	<=	CN_out_sig(3260);
VN_in_sig(3686)	<=	CN_out_sig(3261);
VN_in_sig(4334)	<=	CN_out_sig(3262);
VN_in_sig(4602)	<=	CN_out_sig(3263);
VN_in_sig(238)	<=	CN_out_sig(3264);
VN_in_sig(770)	<=	CN_out_sig(3265);
VN_in_sig(1534)	<=	CN_out_sig(3266);
VN_in_sig(2302)	<=	CN_out_sig(3267);
VN_in_sig(3118)	<=	CN_out_sig(3268);
VN_in_sig(3690)	<=	CN_out_sig(3269);
VN_in_sig(4338)	<=	CN_out_sig(3270);
VN_in_sig(4606)	<=	CN_out_sig(3271);
VN_in_sig(242)	<=	CN_out_sig(3272);
VN_in_sig(774)	<=	CN_out_sig(3273);
VN_in_sig(1538)	<=	CN_out_sig(3274);
VN_in_sig(2306)	<=	CN_out_sig(3275);
VN_in_sig(3122)	<=	CN_out_sig(3276);
VN_in_sig(3694)	<=	CN_out_sig(3277);
VN_in_sig(4342)	<=	CN_out_sig(3278);
VN_in_sig(4610)	<=	CN_out_sig(3279);
VN_in_sig(246)	<=	CN_out_sig(3280);
VN_in_sig(778)	<=	CN_out_sig(3281);
VN_in_sig(1542)	<=	CN_out_sig(3282);
VN_in_sig(2310)	<=	CN_out_sig(3283);
VN_in_sig(3126)	<=	CN_out_sig(3284);
VN_in_sig(3698)	<=	CN_out_sig(3285);
VN_in_sig(4346)	<=	CN_out_sig(3286);
VN_in_sig(4614)	<=	CN_out_sig(3287);
VN_in_sig(250)	<=	CN_out_sig(3288);
VN_in_sig(782)	<=	CN_out_sig(3289);
VN_in_sig(1546)	<=	CN_out_sig(3290);
VN_in_sig(2314)	<=	CN_out_sig(3291);
VN_in_sig(3130)	<=	CN_out_sig(3292);
VN_in_sig(3702)	<=	CN_out_sig(3293);
VN_in_sig(4350)	<=	CN_out_sig(3294);
VN_in_sig(4618)	<=	CN_out_sig(3295);
VN_in_sig(254)	<=	CN_out_sig(3296);
VN_in_sig(786)	<=	CN_out_sig(3297);
VN_in_sig(1550)	<=	CN_out_sig(3298);
VN_in_sig(2318)	<=	CN_out_sig(3299);
VN_in_sig(3134)	<=	CN_out_sig(3300);
VN_in_sig(3706)	<=	CN_out_sig(3301);
VN_in_sig(4354)	<=	CN_out_sig(3302);
VN_in_sig(4622)	<=	CN_out_sig(3303);
VN_in_sig(258)	<=	CN_out_sig(3304);
VN_in_sig(790)	<=	CN_out_sig(3305);
VN_in_sig(1554)	<=	CN_out_sig(3306);
VN_in_sig(2322)	<=	CN_out_sig(3307);
VN_in_sig(3138)	<=	CN_out_sig(3308);
VN_in_sig(3710)	<=	CN_out_sig(3309);
VN_in_sig(4358)	<=	CN_out_sig(3310);
VN_in_sig(4626)	<=	CN_out_sig(3311);
VN_in_sig(262)	<=	CN_out_sig(3312);
VN_in_sig(794)	<=	CN_out_sig(3313);
VN_in_sig(1558)	<=	CN_out_sig(3314);
VN_in_sig(2326)	<=	CN_out_sig(3315);
VN_in_sig(3142)	<=	CN_out_sig(3316);
VN_in_sig(3714)	<=	CN_out_sig(3317);
VN_in_sig(4362)	<=	CN_out_sig(3318);
VN_in_sig(4630)	<=	CN_out_sig(3319);
VN_in_sig(266)	<=	CN_out_sig(3320);
VN_in_sig(798)	<=	CN_out_sig(3321);
VN_in_sig(1562)	<=	CN_out_sig(3322);
VN_in_sig(2330)	<=	CN_out_sig(3323);
VN_in_sig(3146)	<=	CN_out_sig(3324);
VN_in_sig(3718)	<=	CN_out_sig(3325);
VN_in_sig(4366)	<=	CN_out_sig(3326);
VN_in_sig(4634)	<=	CN_out_sig(3327);
VN_in_sig(270)	<=	CN_out_sig(3328);
VN_in_sig(802)	<=	CN_out_sig(3329);
VN_in_sig(1566)	<=	CN_out_sig(3330);
VN_in_sig(2334)	<=	CN_out_sig(3331);
VN_in_sig(3150)	<=	CN_out_sig(3332);
VN_in_sig(3722)	<=	CN_out_sig(3333);
VN_in_sig(4370)	<=	CN_out_sig(3334);
VN_in_sig(4638)	<=	CN_out_sig(3335);
VN_in_sig(274)	<=	CN_out_sig(3336);
VN_in_sig(806)	<=	CN_out_sig(3337);
VN_in_sig(1570)	<=	CN_out_sig(3338);
VN_in_sig(2338)	<=	CN_out_sig(3339);
VN_in_sig(3154)	<=	CN_out_sig(3340);
VN_in_sig(3726)	<=	CN_out_sig(3341);
VN_in_sig(4374)	<=	CN_out_sig(3342);
VN_in_sig(4642)	<=	CN_out_sig(3343);
VN_in_sig(278)	<=	CN_out_sig(3344);
VN_in_sig(810)	<=	CN_out_sig(3345);
VN_in_sig(1574)	<=	CN_out_sig(3346);
VN_in_sig(2342)	<=	CN_out_sig(3347);
VN_in_sig(3158)	<=	CN_out_sig(3348);
VN_in_sig(3730)	<=	CN_out_sig(3349);
VN_in_sig(4378)	<=	CN_out_sig(3350);
VN_in_sig(4646)	<=	CN_out_sig(3351);
VN_in_sig(282)	<=	CN_out_sig(3352);
VN_in_sig(814)	<=	CN_out_sig(3353);
VN_in_sig(1578)	<=	CN_out_sig(3354);
VN_in_sig(2346)	<=	CN_out_sig(3355);
VN_in_sig(3162)	<=	CN_out_sig(3356);
VN_in_sig(3734)	<=	CN_out_sig(3357);
VN_in_sig(4382)	<=	CN_out_sig(3358);
VN_in_sig(4650)	<=	CN_out_sig(3359);
VN_in_sig(286)	<=	CN_out_sig(3360);
VN_in_sig(818)	<=	CN_out_sig(3361);
VN_in_sig(1582)	<=	CN_out_sig(3362);
VN_in_sig(2350)	<=	CN_out_sig(3363);
VN_in_sig(3166)	<=	CN_out_sig(3364);
VN_in_sig(3738)	<=	CN_out_sig(3365);
VN_in_sig(4386)	<=	CN_out_sig(3366);
VN_in_sig(4654)	<=	CN_out_sig(3367);
VN_in_sig(290)	<=	CN_out_sig(3368);
VN_in_sig(822)	<=	CN_out_sig(3369);
VN_in_sig(1586)	<=	CN_out_sig(3370);
VN_in_sig(2354)	<=	CN_out_sig(3371);
VN_in_sig(3170)	<=	CN_out_sig(3372);
VN_in_sig(3742)	<=	CN_out_sig(3373);
VN_in_sig(4390)	<=	CN_out_sig(3374);
VN_in_sig(4658)	<=	CN_out_sig(3375);
VN_in_sig(294)	<=	CN_out_sig(3376);
VN_in_sig(826)	<=	CN_out_sig(3377);
VN_in_sig(1590)	<=	CN_out_sig(3378);
VN_in_sig(2358)	<=	CN_out_sig(3379);
VN_in_sig(3174)	<=	CN_out_sig(3380);
VN_in_sig(3746)	<=	CN_out_sig(3381);
VN_in_sig(4394)	<=	CN_out_sig(3382);
VN_in_sig(4662)	<=	CN_out_sig(3383);
VN_in_sig(298)	<=	CN_out_sig(3384);
VN_in_sig(830)	<=	CN_out_sig(3385);
VN_in_sig(1594)	<=	CN_out_sig(3386);
VN_in_sig(2362)	<=	CN_out_sig(3387);
VN_in_sig(3178)	<=	CN_out_sig(3388);
VN_in_sig(3750)	<=	CN_out_sig(3389);
VN_in_sig(4398)	<=	CN_out_sig(3390);
VN_in_sig(4666)	<=	CN_out_sig(3391);
VN_in_sig(302)	<=	CN_out_sig(3392);
VN_in_sig(834)	<=	CN_out_sig(3393);
VN_in_sig(1598)	<=	CN_out_sig(3394);
VN_in_sig(2366)	<=	CN_out_sig(3395);
VN_in_sig(3182)	<=	CN_out_sig(3396);
VN_in_sig(3754)	<=	CN_out_sig(3397);
VN_in_sig(4402)	<=	CN_out_sig(3398);
VN_in_sig(4670)	<=	CN_out_sig(3399);
VN_in_sig(306)	<=	CN_out_sig(3400);
VN_in_sig(838)	<=	CN_out_sig(3401);
VN_in_sig(1602)	<=	CN_out_sig(3402);
VN_in_sig(2370)	<=	CN_out_sig(3403);
VN_in_sig(3186)	<=	CN_out_sig(3404);
VN_in_sig(3758)	<=	CN_out_sig(3405);
VN_in_sig(4406)	<=	CN_out_sig(3406);
VN_in_sig(4674)	<=	CN_out_sig(3407);
VN_in_sig(310)	<=	CN_out_sig(3408);
VN_in_sig(842)	<=	CN_out_sig(3409);
VN_in_sig(1606)	<=	CN_out_sig(3410);
VN_in_sig(2374)	<=	CN_out_sig(3411);
VN_in_sig(3190)	<=	CN_out_sig(3412);
VN_in_sig(3762)	<=	CN_out_sig(3413);
VN_in_sig(4410)	<=	CN_out_sig(3414);
VN_in_sig(4678)	<=	CN_out_sig(3415);
VN_in_sig(314)	<=	CN_out_sig(3416);
VN_in_sig(846)	<=	CN_out_sig(3417);
VN_in_sig(1610)	<=	CN_out_sig(3418);
VN_in_sig(2162)	<=	CN_out_sig(3419);
VN_in_sig(3194)	<=	CN_out_sig(3420);
VN_in_sig(3766)	<=	CN_out_sig(3421);
VN_in_sig(4414)	<=	CN_out_sig(3422);
VN_in_sig(4682)	<=	CN_out_sig(3423);
VN_in_sig(318)	<=	CN_out_sig(3424);
VN_in_sig(850)	<=	CN_out_sig(3425);
VN_in_sig(1614)	<=	CN_out_sig(3426);
VN_in_sig(2166)	<=	CN_out_sig(3427);
VN_in_sig(3198)	<=	CN_out_sig(3428);
VN_in_sig(3770)	<=	CN_out_sig(3429);
VN_in_sig(4418)	<=	CN_out_sig(3430);
VN_in_sig(4686)	<=	CN_out_sig(3431);
VN_in_sig(322)	<=	CN_out_sig(3432);
VN_in_sig(854)	<=	CN_out_sig(3433);
VN_in_sig(1618)	<=	CN_out_sig(3434);
VN_in_sig(2170)	<=	CN_out_sig(3435);
VN_in_sig(3202)	<=	CN_out_sig(3436);
VN_in_sig(3774)	<=	CN_out_sig(3437);
VN_in_sig(4422)	<=	CN_out_sig(3438);
VN_in_sig(4690)	<=	CN_out_sig(3439);
VN_in_sig(326)	<=	CN_out_sig(3440);
VN_in_sig(858)	<=	CN_out_sig(3441);
VN_in_sig(1622)	<=	CN_out_sig(3442);
VN_in_sig(2174)	<=	CN_out_sig(3443);
VN_in_sig(3206)	<=	CN_out_sig(3444);
VN_in_sig(3778)	<=	CN_out_sig(3445);
VN_in_sig(4426)	<=	CN_out_sig(3446);
VN_in_sig(4694)	<=	CN_out_sig(3447);
VN_in_sig(330)	<=	CN_out_sig(3448);
VN_in_sig(862)	<=	CN_out_sig(3449);
VN_in_sig(1626)	<=	CN_out_sig(3450);
VN_in_sig(2178)	<=	CN_out_sig(3451);
VN_in_sig(3210)	<=	CN_out_sig(3452);
VN_in_sig(3782)	<=	CN_out_sig(3453);
VN_in_sig(4430)	<=	CN_out_sig(3454);
VN_in_sig(4698)	<=	CN_out_sig(3455);
VN_in_sig(38)	<=	CN_out_sig(3456);
VN_in_sig(894)	<=	CN_out_sig(3457);
VN_in_sig(1378)	<=	CN_out_sig(3458);
VN_in_sig(2382)	<=	CN_out_sig(3459);
VN_in_sig(2886)	<=	CN_out_sig(3460);
VN_in_sig(3478)	<=	CN_out_sig(3461);
VN_in_sig(3990)	<=	CN_out_sig(3462);
VN_in_sig(5134)	<=	CN_out_sig(3463);
VN_in_sig(42)	<=	CN_out_sig(3464);
VN_in_sig(898)	<=	CN_out_sig(3465);
VN_in_sig(1382)	<=	CN_out_sig(3466);
VN_in_sig(2386)	<=	CN_out_sig(3467);
VN_in_sig(2890)	<=	CN_out_sig(3468);
VN_in_sig(3482)	<=	CN_out_sig(3469);
VN_in_sig(3994)	<=	CN_out_sig(3470);
VN_in_sig(5138)	<=	CN_out_sig(3471);
VN_in_sig(46)	<=	CN_out_sig(3472);
VN_in_sig(902)	<=	CN_out_sig(3473);
VN_in_sig(1386)	<=	CN_out_sig(3474);
VN_in_sig(2390)	<=	CN_out_sig(3475);
VN_in_sig(2894)	<=	CN_out_sig(3476);
VN_in_sig(3486)	<=	CN_out_sig(3477);
VN_in_sig(3998)	<=	CN_out_sig(3478);
VN_in_sig(5142)	<=	CN_out_sig(3479);
VN_in_sig(50)	<=	CN_out_sig(3480);
VN_in_sig(906)	<=	CN_out_sig(3481);
VN_in_sig(1390)	<=	CN_out_sig(3482);
VN_in_sig(2394)	<=	CN_out_sig(3483);
VN_in_sig(2898)	<=	CN_out_sig(3484);
VN_in_sig(3490)	<=	CN_out_sig(3485);
VN_in_sig(4002)	<=	CN_out_sig(3486);
VN_in_sig(5146)	<=	CN_out_sig(3487);
VN_in_sig(54)	<=	CN_out_sig(3488);
VN_in_sig(910)	<=	CN_out_sig(3489);
VN_in_sig(1394)	<=	CN_out_sig(3490);
VN_in_sig(2398)	<=	CN_out_sig(3491);
VN_in_sig(2902)	<=	CN_out_sig(3492);
VN_in_sig(3494)	<=	CN_out_sig(3493);
VN_in_sig(4006)	<=	CN_out_sig(3494);
VN_in_sig(5150)	<=	CN_out_sig(3495);
VN_in_sig(58)	<=	CN_out_sig(3496);
VN_in_sig(914)	<=	CN_out_sig(3497);
VN_in_sig(1398)	<=	CN_out_sig(3498);
VN_in_sig(2402)	<=	CN_out_sig(3499);
VN_in_sig(2906)	<=	CN_out_sig(3500);
VN_in_sig(3498)	<=	CN_out_sig(3501);
VN_in_sig(4010)	<=	CN_out_sig(3502);
VN_in_sig(5154)	<=	CN_out_sig(3503);
VN_in_sig(62)	<=	CN_out_sig(3504);
VN_in_sig(918)	<=	CN_out_sig(3505);
VN_in_sig(1402)	<=	CN_out_sig(3506);
VN_in_sig(2406)	<=	CN_out_sig(3507);
VN_in_sig(2910)	<=	CN_out_sig(3508);
VN_in_sig(3502)	<=	CN_out_sig(3509);
VN_in_sig(4014)	<=	CN_out_sig(3510);
VN_in_sig(5158)	<=	CN_out_sig(3511);
VN_in_sig(66)	<=	CN_out_sig(3512);
VN_in_sig(922)	<=	CN_out_sig(3513);
VN_in_sig(1406)	<=	CN_out_sig(3514);
VN_in_sig(2410)	<=	CN_out_sig(3515);
VN_in_sig(2914)	<=	CN_out_sig(3516);
VN_in_sig(3506)	<=	CN_out_sig(3517);
VN_in_sig(4018)	<=	CN_out_sig(3518);
VN_in_sig(5162)	<=	CN_out_sig(3519);
VN_in_sig(70)	<=	CN_out_sig(3520);
VN_in_sig(926)	<=	CN_out_sig(3521);
VN_in_sig(1410)	<=	CN_out_sig(3522);
VN_in_sig(2414)	<=	CN_out_sig(3523);
VN_in_sig(2918)	<=	CN_out_sig(3524);
VN_in_sig(3510)	<=	CN_out_sig(3525);
VN_in_sig(4022)	<=	CN_out_sig(3526);
VN_in_sig(5166)	<=	CN_out_sig(3527);
VN_in_sig(74)	<=	CN_out_sig(3528);
VN_in_sig(930)	<=	CN_out_sig(3529);
VN_in_sig(1414)	<=	CN_out_sig(3530);
VN_in_sig(2418)	<=	CN_out_sig(3531);
VN_in_sig(2922)	<=	CN_out_sig(3532);
VN_in_sig(3514)	<=	CN_out_sig(3533);
VN_in_sig(4026)	<=	CN_out_sig(3534);
VN_in_sig(5170)	<=	CN_out_sig(3535);
VN_in_sig(78)	<=	CN_out_sig(3536);
VN_in_sig(934)	<=	CN_out_sig(3537);
VN_in_sig(1418)	<=	CN_out_sig(3538);
VN_in_sig(2422)	<=	CN_out_sig(3539);
VN_in_sig(2926)	<=	CN_out_sig(3540);
VN_in_sig(3518)	<=	CN_out_sig(3541);
VN_in_sig(4030)	<=	CN_out_sig(3542);
VN_in_sig(5174)	<=	CN_out_sig(3543);
VN_in_sig(82)	<=	CN_out_sig(3544);
VN_in_sig(938)	<=	CN_out_sig(3545);
VN_in_sig(1422)	<=	CN_out_sig(3546);
VN_in_sig(2426)	<=	CN_out_sig(3547);
VN_in_sig(2930)	<=	CN_out_sig(3548);
VN_in_sig(3522)	<=	CN_out_sig(3549);
VN_in_sig(4034)	<=	CN_out_sig(3550);
VN_in_sig(5178)	<=	CN_out_sig(3551);
VN_in_sig(86)	<=	CN_out_sig(3552);
VN_in_sig(942)	<=	CN_out_sig(3553);
VN_in_sig(1426)	<=	CN_out_sig(3554);
VN_in_sig(2430)	<=	CN_out_sig(3555);
VN_in_sig(2934)	<=	CN_out_sig(3556);
VN_in_sig(3526)	<=	CN_out_sig(3557);
VN_in_sig(4038)	<=	CN_out_sig(3558);
VN_in_sig(5182)	<=	CN_out_sig(3559);
VN_in_sig(90)	<=	CN_out_sig(3560);
VN_in_sig(946)	<=	CN_out_sig(3561);
VN_in_sig(1430)	<=	CN_out_sig(3562);
VN_in_sig(2434)	<=	CN_out_sig(3563);
VN_in_sig(2938)	<=	CN_out_sig(3564);
VN_in_sig(3530)	<=	CN_out_sig(3565);
VN_in_sig(4042)	<=	CN_out_sig(3566);
VN_in_sig(4970)	<=	CN_out_sig(3567);
VN_in_sig(94)	<=	CN_out_sig(3568);
VN_in_sig(950)	<=	CN_out_sig(3569);
VN_in_sig(1434)	<=	CN_out_sig(3570);
VN_in_sig(2438)	<=	CN_out_sig(3571);
VN_in_sig(2942)	<=	CN_out_sig(3572);
VN_in_sig(3534)	<=	CN_out_sig(3573);
VN_in_sig(4046)	<=	CN_out_sig(3574);
VN_in_sig(4974)	<=	CN_out_sig(3575);
VN_in_sig(98)	<=	CN_out_sig(3576);
VN_in_sig(954)	<=	CN_out_sig(3577);
VN_in_sig(1438)	<=	CN_out_sig(3578);
VN_in_sig(2442)	<=	CN_out_sig(3579);
VN_in_sig(2946)	<=	CN_out_sig(3580);
VN_in_sig(3538)	<=	CN_out_sig(3581);
VN_in_sig(4050)	<=	CN_out_sig(3582);
VN_in_sig(4978)	<=	CN_out_sig(3583);
VN_in_sig(102)	<=	CN_out_sig(3584);
VN_in_sig(958)	<=	CN_out_sig(3585);
VN_in_sig(1442)	<=	CN_out_sig(3586);
VN_in_sig(2446)	<=	CN_out_sig(3587);
VN_in_sig(2950)	<=	CN_out_sig(3588);
VN_in_sig(3542)	<=	CN_out_sig(3589);
VN_in_sig(4054)	<=	CN_out_sig(3590);
VN_in_sig(4982)	<=	CN_out_sig(3591);
VN_in_sig(106)	<=	CN_out_sig(3592);
VN_in_sig(962)	<=	CN_out_sig(3593);
VN_in_sig(1446)	<=	CN_out_sig(3594);
VN_in_sig(2450)	<=	CN_out_sig(3595);
VN_in_sig(2954)	<=	CN_out_sig(3596);
VN_in_sig(3546)	<=	CN_out_sig(3597);
VN_in_sig(4058)	<=	CN_out_sig(3598);
VN_in_sig(4986)	<=	CN_out_sig(3599);
VN_in_sig(110)	<=	CN_out_sig(3600);
VN_in_sig(966)	<=	CN_out_sig(3601);
VN_in_sig(1450)	<=	CN_out_sig(3602);
VN_in_sig(2454)	<=	CN_out_sig(3603);
VN_in_sig(2958)	<=	CN_out_sig(3604);
VN_in_sig(3550)	<=	CN_out_sig(3605);
VN_in_sig(4062)	<=	CN_out_sig(3606);
VN_in_sig(4990)	<=	CN_out_sig(3607);
VN_in_sig(114)	<=	CN_out_sig(3608);
VN_in_sig(970)	<=	CN_out_sig(3609);
VN_in_sig(1454)	<=	CN_out_sig(3610);
VN_in_sig(2458)	<=	CN_out_sig(3611);
VN_in_sig(2962)	<=	CN_out_sig(3612);
VN_in_sig(3554)	<=	CN_out_sig(3613);
VN_in_sig(4066)	<=	CN_out_sig(3614);
VN_in_sig(4994)	<=	CN_out_sig(3615);
VN_in_sig(118)	<=	CN_out_sig(3616);
VN_in_sig(974)	<=	CN_out_sig(3617);
VN_in_sig(1458)	<=	CN_out_sig(3618);
VN_in_sig(2462)	<=	CN_out_sig(3619);
VN_in_sig(2966)	<=	CN_out_sig(3620);
VN_in_sig(3558)	<=	CN_out_sig(3621);
VN_in_sig(4070)	<=	CN_out_sig(3622);
VN_in_sig(4998)	<=	CN_out_sig(3623);
VN_in_sig(122)	<=	CN_out_sig(3624);
VN_in_sig(978)	<=	CN_out_sig(3625);
VN_in_sig(1462)	<=	CN_out_sig(3626);
VN_in_sig(2466)	<=	CN_out_sig(3627);
VN_in_sig(2970)	<=	CN_out_sig(3628);
VN_in_sig(3562)	<=	CN_out_sig(3629);
VN_in_sig(4074)	<=	CN_out_sig(3630);
VN_in_sig(5002)	<=	CN_out_sig(3631);
VN_in_sig(126)	<=	CN_out_sig(3632);
VN_in_sig(982)	<=	CN_out_sig(3633);
VN_in_sig(1466)	<=	CN_out_sig(3634);
VN_in_sig(2470)	<=	CN_out_sig(3635);
VN_in_sig(2974)	<=	CN_out_sig(3636);
VN_in_sig(3566)	<=	CN_out_sig(3637);
VN_in_sig(4078)	<=	CN_out_sig(3638);
VN_in_sig(5006)	<=	CN_out_sig(3639);
VN_in_sig(130)	<=	CN_out_sig(3640);
VN_in_sig(986)	<=	CN_out_sig(3641);
VN_in_sig(1470)	<=	CN_out_sig(3642);
VN_in_sig(2474)	<=	CN_out_sig(3643);
VN_in_sig(2978)	<=	CN_out_sig(3644);
VN_in_sig(3570)	<=	CN_out_sig(3645);
VN_in_sig(4082)	<=	CN_out_sig(3646);
VN_in_sig(5010)	<=	CN_out_sig(3647);
VN_in_sig(134)	<=	CN_out_sig(3648);
VN_in_sig(990)	<=	CN_out_sig(3649);
VN_in_sig(1474)	<=	CN_out_sig(3650);
VN_in_sig(2478)	<=	CN_out_sig(3651);
VN_in_sig(2982)	<=	CN_out_sig(3652);
VN_in_sig(3574)	<=	CN_out_sig(3653);
VN_in_sig(4086)	<=	CN_out_sig(3654);
VN_in_sig(5014)	<=	CN_out_sig(3655);
VN_in_sig(138)	<=	CN_out_sig(3656);
VN_in_sig(994)	<=	CN_out_sig(3657);
VN_in_sig(1478)	<=	CN_out_sig(3658);
VN_in_sig(2482)	<=	CN_out_sig(3659);
VN_in_sig(2986)	<=	CN_out_sig(3660);
VN_in_sig(3578)	<=	CN_out_sig(3661);
VN_in_sig(4090)	<=	CN_out_sig(3662);
VN_in_sig(5018)	<=	CN_out_sig(3663);
VN_in_sig(142)	<=	CN_out_sig(3664);
VN_in_sig(998)	<=	CN_out_sig(3665);
VN_in_sig(1482)	<=	CN_out_sig(3666);
VN_in_sig(2486)	<=	CN_out_sig(3667);
VN_in_sig(2990)	<=	CN_out_sig(3668);
VN_in_sig(3582)	<=	CN_out_sig(3669);
VN_in_sig(4094)	<=	CN_out_sig(3670);
VN_in_sig(5022)	<=	CN_out_sig(3671);
VN_in_sig(146)	<=	CN_out_sig(3672);
VN_in_sig(1002)	<=	CN_out_sig(3673);
VN_in_sig(1486)	<=	CN_out_sig(3674);
VN_in_sig(2490)	<=	CN_out_sig(3675);
VN_in_sig(2994)	<=	CN_out_sig(3676);
VN_in_sig(3586)	<=	CN_out_sig(3677);
VN_in_sig(4098)	<=	CN_out_sig(3678);
VN_in_sig(5026)	<=	CN_out_sig(3679);
VN_in_sig(150)	<=	CN_out_sig(3680);
VN_in_sig(1006)	<=	CN_out_sig(3681);
VN_in_sig(1490)	<=	CN_out_sig(3682);
VN_in_sig(2494)	<=	CN_out_sig(3683);
VN_in_sig(2998)	<=	CN_out_sig(3684);
VN_in_sig(3590)	<=	CN_out_sig(3685);
VN_in_sig(4102)	<=	CN_out_sig(3686);
VN_in_sig(5030)	<=	CN_out_sig(3687);
VN_in_sig(154)	<=	CN_out_sig(3688);
VN_in_sig(1010)	<=	CN_out_sig(3689);
VN_in_sig(1494)	<=	CN_out_sig(3690);
VN_in_sig(2498)	<=	CN_out_sig(3691);
VN_in_sig(3002)	<=	CN_out_sig(3692);
VN_in_sig(3594)	<=	CN_out_sig(3693);
VN_in_sig(3890)	<=	CN_out_sig(3694);
VN_in_sig(5034)	<=	CN_out_sig(3695);
VN_in_sig(158)	<=	CN_out_sig(3696);
VN_in_sig(1014)	<=	CN_out_sig(3697);
VN_in_sig(1498)	<=	CN_out_sig(3698);
VN_in_sig(2502)	<=	CN_out_sig(3699);
VN_in_sig(3006)	<=	CN_out_sig(3700);
VN_in_sig(3598)	<=	CN_out_sig(3701);
VN_in_sig(3894)	<=	CN_out_sig(3702);
VN_in_sig(5038)	<=	CN_out_sig(3703);
VN_in_sig(162)	<=	CN_out_sig(3704);
VN_in_sig(1018)	<=	CN_out_sig(3705);
VN_in_sig(1502)	<=	CN_out_sig(3706);
VN_in_sig(2506)	<=	CN_out_sig(3707);
VN_in_sig(3010)	<=	CN_out_sig(3708);
VN_in_sig(3602)	<=	CN_out_sig(3709);
VN_in_sig(3898)	<=	CN_out_sig(3710);
VN_in_sig(5042)	<=	CN_out_sig(3711);
VN_in_sig(166)	<=	CN_out_sig(3712);
VN_in_sig(1022)	<=	CN_out_sig(3713);
VN_in_sig(1506)	<=	CN_out_sig(3714);
VN_in_sig(2510)	<=	CN_out_sig(3715);
VN_in_sig(3014)	<=	CN_out_sig(3716);
VN_in_sig(3606)	<=	CN_out_sig(3717);
VN_in_sig(3902)	<=	CN_out_sig(3718);
VN_in_sig(5046)	<=	CN_out_sig(3719);
VN_in_sig(170)	<=	CN_out_sig(3720);
VN_in_sig(1026)	<=	CN_out_sig(3721);
VN_in_sig(1510)	<=	CN_out_sig(3722);
VN_in_sig(2514)	<=	CN_out_sig(3723);
VN_in_sig(3018)	<=	CN_out_sig(3724);
VN_in_sig(3610)	<=	CN_out_sig(3725);
VN_in_sig(3906)	<=	CN_out_sig(3726);
VN_in_sig(5050)	<=	CN_out_sig(3727);
VN_in_sig(174)	<=	CN_out_sig(3728);
VN_in_sig(1030)	<=	CN_out_sig(3729);
VN_in_sig(1298)	<=	CN_out_sig(3730);
VN_in_sig(2518)	<=	CN_out_sig(3731);
VN_in_sig(3022)	<=	CN_out_sig(3732);
VN_in_sig(3614)	<=	CN_out_sig(3733);
VN_in_sig(3910)	<=	CN_out_sig(3734);
VN_in_sig(5054)	<=	CN_out_sig(3735);
VN_in_sig(178)	<=	CN_out_sig(3736);
VN_in_sig(1034)	<=	CN_out_sig(3737);
VN_in_sig(1302)	<=	CN_out_sig(3738);
VN_in_sig(2522)	<=	CN_out_sig(3739);
VN_in_sig(2810)	<=	CN_out_sig(3740);
VN_in_sig(3618)	<=	CN_out_sig(3741);
VN_in_sig(3914)	<=	CN_out_sig(3742);
VN_in_sig(5058)	<=	CN_out_sig(3743);
VN_in_sig(182)	<=	CN_out_sig(3744);
VN_in_sig(1038)	<=	CN_out_sig(3745);
VN_in_sig(1306)	<=	CN_out_sig(3746);
VN_in_sig(2526)	<=	CN_out_sig(3747);
VN_in_sig(2814)	<=	CN_out_sig(3748);
VN_in_sig(3622)	<=	CN_out_sig(3749);
VN_in_sig(3918)	<=	CN_out_sig(3750);
VN_in_sig(5062)	<=	CN_out_sig(3751);
VN_in_sig(186)	<=	CN_out_sig(3752);
VN_in_sig(1042)	<=	CN_out_sig(3753);
VN_in_sig(1310)	<=	CN_out_sig(3754);
VN_in_sig(2530)	<=	CN_out_sig(3755);
VN_in_sig(2818)	<=	CN_out_sig(3756);
VN_in_sig(3626)	<=	CN_out_sig(3757);
VN_in_sig(3922)	<=	CN_out_sig(3758);
VN_in_sig(5066)	<=	CN_out_sig(3759);
VN_in_sig(190)	<=	CN_out_sig(3760);
VN_in_sig(1046)	<=	CN_out_sig(3761);
VN_in_sig(1314)	<=	CN_out_sig(3762);
VN_in_sig(2534)	<=	CN_out_sig(3763);
VN_in_sig(2822)	<=	CN_out_sig(3764);
VN_in_sig(3630)	<=	CN_out_sig(3765);
VN_in_sig(3926)	<=	CN_out_sig(3766);
VN_in_sig(5070)	<=	CN_out_sig(3767);
VN_in_sig(194)	<=	CN_out_sig(3768);
VN_in_sig(1050)	<=	CN_out_sig(3769);
VN_in_sig(1318)	<=	CN_out_sig(3770);
VN_in_sig(2538)	<=	CN_out_sig(3771);
VN_in_sig(2826)	<=	CN_out_sig(3772);
VN_in_sig(3634)	<=	CN_out_sig(3773);
VN_in_sig(3930)	<=	CN_out_sig(3774);
VN_in_sig(5074)	<=	CN_out_sig(3775);
VN_in_sig(198)	<=	CN_out_sig(3776);
VN_in_sig(1054)	<=	CN_out_sig(3777);
VN_in_sig(1322)	<=	CN_out_sig(3778);
VN_in_sig(2542)	<=	CN_out_sig(3779);
VN_in_sig(2830)	<=	CN_out_sig(3780);
VN_in_sig(3638)	<=	CN_out_sig(3781);
VN_in_sig(3934)	<=	CN_out_sig(3782);
VN_in_sig(5078)	<=	CN_out_sig(3783);
VN_in_sig(202)	<=	CN_out_sig(3784);
VN_in_sig(1058)	<=	CN_out_sig(3785);
VN_in_sig(1326)	<=	CN_out_sig(3786);
VN_in_sig(2546)	<=	CN_out_sig(3787);
VN_in_sig(2834)	<=	CN_out_sig(3788);
VN_in_sig(3642)	<=	CN_out_sig(3789);
VN_in_sig(3938)	<=	CN_out_sig(3790);
VN_in_sig(5082)	<=	CN_out_sig(3791);
VN_in_sig(206)	<=	CN_out_sig(3792);
VN_in_sig(1062)	<=	CN_out_sig(3793);
VN_in_sig(1330)	<=	CN_out_sig(3794);
VN_in_sig(2550)	<=	CN_out_sig(3795);
VN_in_sig(2838)	<=	CN_out_sig(3796);
VN_in_sig(3646)	<=	CN_out_sig(3797);
VN_in_sig(3942)	<=	CN_out_sig(3798);
VN_in_sig(5086)	<=	CN_out_sig(3799);
VN_in_sig(210)	<=	CN_out_sig(3800);
VN_in_sig(1066)	<=	CN_out_sig(3801);
VN_in_sig(1334)	<=	CN_out_sig(3802);
VN_in_sig(2554)	<=	CN_out_sig(3803);
VN_in_sig(2842)	<=	CN_out_sig(3804);
VN_in_sig(3650)	<=	CN_out_sig(3805);
VN_in_sig(3946)	<=	CN_out_sig(3806);
VN_in_sig(5090)	<=	CN_out_sig(3807);
VN_in_sig(214)	<=	CN_out_sig(3808);
VN_in_sig(1070)	<=	CN_out_sig(3809);
VN_in_sig(1338)	<=	CN_out_sig(3810);
VN_in_sig(2558)	<=	CN_out_sig(3811);
VN_in_sig(2846)	<=	CN_out_sig(3812);
VN_in_sig(3654)	<=	CN_out_sig(3813);
VN_in_sig(3950)	<=	CN_out_sig(3814);
VN_in_sig(5094)	<=	CN_out_sig(3815);
VN_in_sig(2)	<=	CN_out_sig(3816);
VN_in_sig(1074)	<=	CN_out_sig(3817);
VN_in_sig(1342)	<=	CN_out_sig(3818);
VN_in_sig(2562)	<=	CN_out_sig(3819);
VN_in_sig(2850)	<=	CN_out_sig(3820);
VN_in_sig(3658)	<=	CN_out_sig(3821);
VN_in_sig(3954)	<=	CN_out_sig(3822);
VN_in_sig(5098)	<=	CN_out_sig(3823);
VN_in_sig(6)	<=	CN_out_sig(3824);
VN_in_sig(1078)	<=	CN_out_sig(3825);
VN_in_sig(1346)	<=	CN_out_sig(3826);
VN_in_sig(2566)	<=	CN_out_sig(3827);
VN_in_sig(2854)	<=	CN_out_sig(3828);
VN_in_sig(3662)	<=	CN_out_sig(3829);
VN_in_sig(3958)	<=	CN_out_sig(3830);
VN_in_sig(5102)	<=	CN_out_sig(3831);
VN_in_sig(10)	<=	CN_out_sig(3832);
VN_in_sig(866)	<=	CN_out_sig(3833);
VN_in_sig(1350)	<=	CN_out_sig(3834);
VN_in_sig(2570)	<=	CN_out_sig(3835);
VN_in_sig(2858)	<=	CN_out_sig(3836);
VN_in_sig(3666)	<=	CN_out_sig(3837);
VN_in_sig(3962)	<=	CN_out_sig(3838);
VN_in_sig(5106)	<=	CN_out_sig(3839);
VN_in_sig(14)	<=	CN_out_sig(3840);
VN_in_sig(870)	<=	CN_out_sig(3841);
VN_in_sig(1354)	<=	CN_out_sig(3842);
VN_in_sig(2574)	<=	CN_out_sig(3843);
VN_in_sig(2862)	<=	CN_out_sig(3844);
VN_in_sig(3670)	<=	CN_out_sig(3845);
VN_in_sig(3966)	<=	CN_out_sig(3846);
VN_in_sig(5110)	<=	CN_out_sig(3847);
VN_in_sig(18)	<=	CN_out_sig(3848);
VN_in_sig(874)	<=	CN_out_sig(3849);
VN_in_sig(1358)	<=	CN_out_sig(3850);
VN_in_sig(2578)	<=	CN_out_sig(3851);
VN_in_sig(2866)	<=	CN_out_sig(3852);
VN_in_sig(3458)	<=	CN_out_sig(3853);
VN_in_sig(3970)	<=	CN_out_sig(3854);
VN_in_sig(5114)	<=	CN_out_sig(3855);
VN_in_sig(22)	<=	CN_out_sig(3856);
VN_in_sig(878)	<=	CN_out_sig(3857);
VN_in_sig(1362)	<=	CN_out_sig(3858);
VN_in_sig(2582)	<=	CN_out_sig(3859);
VN_in_sig(2870)	<=	CN_out_sig(3860);
VN_in_sig(3462)	<=	CN_out_sig(3861);
VN_in_sig(3974)	<=	CN_out_sig(3862);
VN_in_sig(5118)	<=	CN_out_sig(3863);
VN_in_sig(26)	<=	CN_out_sig(3864);
VN_in_sig(882)	<=	CN_out_sig(3865);
VN_in_sig(1366)	<=	CN_out_sig(3866);
VN_in_sig(2586)	<=	CN_out_sig(3867);
VN_in_sig(2874)	<=	CN_out_sig(3868);
VN_in_sig(3466)	<=	CN_out_sig(3869);
VN_in_sig(3978)	<=	CN_out_sig(3870);
VN_in_sig(5122)	<=	CN_out_sig(3871);
VN_in_sig(30)	<=	CN_out_sig(3872);
VN_in_sig(886)	<=	CN_out_sig(3873);
VN_in_sig(1370)	<=	CN_out_sig(3874);
VN_in_sig(2590)	<=	CN_out_sig(3875);
VN_in_sig(2878)	<=	CN_out_sig(3876);
VN_in_sig(3470)	<=	CN_out_sig(3877);
VN_in_sig(3982)	<=	CN_out_sig(3878);
VN_in_sig(5126)	<=	CN_out_sig(3879);
VN_in_sig(34)	<=	CN_out_sig(3880);
VN_in_sig(890)	<=	CN_out_sig(3881);
VN_in_sig(1374)	<=	CN_out_sig(3882);
VN_in_sig(2378)	<=	CN_out_sig(3883);
VN_in_sig(2882)	<=	CN_out_sig(3884);
VN_in_sig(3474)	<=	CN_out_sig(3885);
VN_in_sig(3986)	<=	CN_out_sig(3886);
VN_in_sig(5130)	<=	CN_out_sig(3887);
VN_in_sig(647)	<=	CN_out_sig(3888);
VN_in_sig(1095)	<=	CN_out_sig(3889);
VN_in_sig(1835)	<=	CN_out_sig(3890);
VN_in_sig(2175)	<=	CN_out_sig(3891);
VN_in_sig(3147)	<=	CN_out_sig(3892);
VN_in_sig(3695)	<=	CN_out_sig(3893);
VN_in_sig(4247)	<=	CN_out_sig(3894);
VN_in_sig(4931)	<=	CN_out_sig(3895);
VN_in_sig(435)	<=	CN_out_sig(3896);
VN_in_sig(1099)	<=	CN_out_sig(3897);
VN_in_sig(1839)	<=	CN_out_sig(3898);
VN_in_sig(2179)	<=	CN_out_sig(3899);
VN_in_sig(3151)	<=	CN_out_sig(3900);
VN_in_sig(3699)	<=	CN_out_sig(3901);
VN_in_sig(4251)	<=	CN_out_sig(3902);
VN_in_sig(4935)	<=	CN_out_sig(3903);
VN_in_sig(439)	<=	CN_out_sig(3904);
VN_in_sig(1103)	<=	CN_out_sig(3905);
VN_in_sig(1843)	<=	CN_out_sig(3906);
VN_in_sig(2183)	<=	CN_out_sig(3907);
VN_in_sig(3155)	<=	CN_out_sig(3908);
VN_in_sig(3703)	<=	CN_out_sig(3909);
VN_in_sig(4255)	<=	CN_out_sig(3910);
VN_in_sig(4939)	<=	CN_out_sig(3911);
VN_in_sig(443)	<=	CN_out_sig(3912);
VN_in_sig(1107)	<=	CN_out_sig(3913);
VN_in_sig(1847)	<=	CN_out_sig(3914);
VN_in_sig(2187)	<=	CN_out_sig(3915);
VN_in_sig(3159)	<=	CN_out_sig(3916);
VN_in_sig(3707)	<=	CN_out_sig(3917);
VN_in_sig(4259)	<=	CN_out_sig(3918);
VN_in_sig(4943)	<=	CN_out_sig(3919);
VN_in_sig(447)	<=	CN_out_sig(3920);
VN_in_sig(1111)	<=	CN_out_sig(3921);
VN_in_sig(1851)	<=	CN_out_sig(3922);
VN_in_sig(2191)	<=	CN_out_sig(3923);
VN_in_sig(3163)	<=	CN_out_sig(3924);
VN_in_sig(3711)	<=	CN_out_sig(3925);
VN_in_sig(4263)	<=	CN_out_sig(3926);
VN_in_sig(4947)	<=	CN_out_sig(3927);
VN_in_sig(451)	<=	CN_out_sig(3928);
VN_in_sig(1115)	<=	CN_out_sig(3929);
VN_in_sig(1855)	<=	CN_out_sig(3930);
VN_in_sig(2195)	<=	CN_out_sig(3931);
VN_in_sig(3167)	<=	CN_out_sig(3932);
VN_in_sig(3715)	<=	CN_out_sig(3933);
VN_in_sig(4267)	<=	CN_out_sig(3934);
VN_in_sig(4951)	<=	CN_out_sig(3935);
VN_in_sig(455)	<=	CN_out_sig(3936);
VN_in_sig(1119)	<=	CN_out_sig(3937);
VN_in_sig(1859)	<=	CN_out_sig(3938);
VN_in_sig(2199)	<=	CN_out_sig(3939);
VN_in_sig(3171)	<=	CN_out_sig(3940);
VN_in_sig(3719)	<=	CN_out_sig(3941);
VN_in_sig(4271)	<=	CN_out_sig(3942);
VN_in_sig(4955)	<=	CN_out_sig(3943);
VN_in_sig(459)	<=	CN_out_sig(3944);
VN_in_sig(1123)	<=	CN_out_sig(3945);
VN_in_sig(1863)	<=	CN_out_sig(3946);
VN_in_sig(2203)	<=	CN_out_sig(3947);
VN_in_sig(3175)	<=	CN_out_sig(3948);
VN_in_sig(3723)	<=	CN_out_sig(3949);
VN_in_sig(4275)	<=	CN_out_sig(3950);
VN_in_sig(4959)	<=	CN_out_sig(3951);
VN_in_sig(463)	<=	CN_out_sig(3952);
VN_in_sig(1127)	<=	CN_out_sig(3953);
VN_in_sig(1867)	<=	CN_out_sig(3954);
VN_in_sig(2207)	<=	CN_out_sig(3955);
VN_in_sig(3179)	<=	CN_out_sig(3956);
VN_in_sig(3727)	<=	CN_out_sig(3957);
VN_in_sig(4279)	<=	CN_out_sig(3958);
VN_in_sig(4963)	<=	CN_out_sig(3959);
VN_in_sig(467)	<=	CN_out_sig(3960);
VN_in_sig(1131)	<=	CN_out_sig(3961);
VN_in_sig(1871)	<=	CN_out_sig(3962);
VN_in_sig(2211)	<=	CN_out_sig(3963);
VN_in_sig(3183)	<=	CN_out_sig(3964);
VN_in_sig(3731)	<=	CN_out_sig(3965);
VN_in_sig(4283)	<=	CN_out_sig(3966);
VN_in_sig(4967)	<=	CN_out_sig(3967);
VN_in_sig(471)	<=	CN_out_sig(3968);
VN_in_sig(1135)	<=	CN_out_sig(3969);
VN_in_sig(1875)	<=	CN_out_sig(3970);
VN_in_sig(2215)	<=	CN_out_sig(3971);
VN_in_sig(3187)	<=	CN_out_sig(3972);
VN_in_sig(3735)	<=	CN_out_sig(3973);
VN_in_sig(4287)	<=	CN_out_sig(3974);
VN_in_sig(4755)	<=	CN_out_sig(3975);
VN_in_sig(475)	<=	CN_out_sig(3976);
VN_in_sig(1139)	<=	CN_out_sig(3977);
VN_in_sig(1879)	<=	CN_out_sig(3978);
VN_in_sig(2219)	<=	CN_out_sig(3979);
VN_in_sig(3191)	<=	CN_out_sig(3980);
VN_in_sig(3739)	<=	CN_out_sig(3981);
VN_in_sig(4291)	<=	CN_out_sig(3982);
VN_in_sig(4759)	<=	CN_out_sig(3983);
VN_in_sig(479)	<=	CN_out_sig(3984);
VN_in_sig(1143)	<=	CN_out_sig(3985);
VN_in_sig(1883)	<=	CN_out_sig(3986);
VN_in_sig(2223)	<=	CN_out_sig(3987);
VN_in_sig(3195)	<=	CN_out_sig(3988);
VN_in_sig(3743)	<=	CN_out_sig(3989);
VN_in_sig(4295)	<=	CN_out_sig(3990);
VN_in_sig(4763)	<=	CN_out_sig(3991);
VN_in_sig(483)	<=	CN_out_sig(3992);
VN_in_sig(1147)	<=	CN_out_sig(3993);
VN_in_sig(1887)	<=	CN_out_sig(3994);
VN_in_sig(2227)	<=	CN_out_sig(3995);
VN_in_sig(3199)	<=	CN_out_sig(3996);
VN_in_sig(3747)	<=	CN_out_sig(3997);
VN_in_sig(4299)	<=	CN_out_sig(3998);
VN_in_sig(4767)	<=	CN_out_sig(3999);
VN_in_sig(487)	<=	CN_out_sig(4000);
VN_in_sig(1151)	<=	CN_out_sig(4001);
VN_in_sig(1891)	<=	CN_out_sig(4002);
VN_in_sig(2231)	<=	CN_out_sig(4003);
VN_in_sig(3203)	<=	CN_out_sig(4004);
VN_in_sig(3751)	<=	CN_out_sig(4005);
VN_in_sig(4303)	<=	CN_out_sig(4006);
VN_in_sig(4771)	<=	CN_out_sig(4007);
VN_in_sig(491)	<=	CN_out_sig(4008);
VN_in_sig(1155)	<=	CN_out_sig(4009);
VN_in_sig(1895)	<=	CN_out_sig(4010);
VN_in_sig(2235)	<=	CN_out_sig(4011);
VN_in_sig(3207)	<=	CN_out_sig(4012);
VN_in_sig(3755)	<=	CN_out_sig(4013);
VN_in_sig(4307)	<=	CN_out_sig(4014);
VN_in_sig(4775)	<=	CN_out_sig(4015);
VN_in_sig(495)	<=	CN_out_sig(4016);
VN_in_sig(1159)	<=	CN_out_sig(4017);
VN_in_sig(1899)	<=	CN_out_sig(4018);
VN_in_sig(2239)	<=	CN_out_sig(4019);
VN_in_sig(3211)	<=	CN_out_sig(4020);
VN_in_sig(3759)	<=	CN_out_sig(4021);
VN_in_sig(4311)	<=	CN_out_sig(4022);
VN_in_sig(4779)	<=	CN_out_sig(4023);
VN_in_sig(499)	<=	CN_out_sig(4024);
VN_in_sig(1163)	<=	CN_out_sig(4025);
VN_in_sig(1903)	<=	CN_out_sig(4026);
VN_in_sig(2243)	<=	CN_out_sig(4027);
VN_in_sig(3215)	<=	CN_out_sig(4028);
VN_in_sig(3763)	<=	CN_out_sig(4029);
VN_in_sig(4315)	<=	CN_out_sig(4030);
VN_in_sig(4783)	<=	CN_out_sig(4031);
VN_in_sig(503)	<=	CN_out_sig(4032);
VN_in_sig(1167)	<=	CN_out_sig(4033);
VN_in_sig(1907)	<=	CN_out_sig(4034);
VN_in_sig(2247)	<=	CN_out_sig(4035);
VN_in_sig(3219)	<=	CN_out_sig(4036);
VN_in_sig(3767)	<=	CN_out_sig(4037);
VN_in_sig(4319)	<=	CN_out_sig(4038);
VN_in_sig(4787)	<=	CN_out_sig(4039);
VN_in_sig(507)	<=	CN_out_sig(4040);
VN_in_sig(1171)	<=	CN_out_sig(4041);
VN_in_sig(1911)	<=	CN_out_sig(4042);
VN_in_sig(2251)	<=	CN_out_sig(4043);
VN_in_sig(3223)	<=	CN_out_sig(4044);
VN_in_sig(3771)	<=	CN_out_sig(4045);
VN_in_sig(4107)	<=	CN_out_sig(4046);
VN_in_sig(4791)	<=	CN_out_sig(4047);
VN_in_sig(511)	<=	CN_out_sig(4048);
VN_in_sig(1175)	<=	CN_out_sig(4049);
VN_in_sig(1915)	<=	CN_out_sig(4050);
VN_in_sig(2255)	<=	CN_out_sig(4051);
VN_in_sig(3227)	<=	CN_out_sig(4052);
VN_in_sig(3775)	<=	CN_out_sig(4053);
VN_in_sig(4111)	<=	CN_out_sig(4054);
VN_in_sig(4795)	<=	CN_out_sig(4055);
VN_in_sig(515)	<=	CN_out_sig(4056);
VN_in_sig(1179)	<=	CN_out_sig(4057);
VN_in_sig(1919)	<=	CN_out_sig(4058);
VN_in_sig(2259)	<=	CN_out_sig(4059);
VN_in_sig(3231)	<=	CN_out_sig(4060);
VN_in_sig(3779)	<=	CN_out_sig(4061);
VN_in_sig(4115)	<=	CN_out_sig(4062);
VN_in_sig(4799)	<=	CN_out_sig(4063);
VN_in_sig(519)	<=	CN_out_sig(4064);
VN_in_sig(1183)	<=	CN_out_sig(4065);
VN_in_sig(1923)	<=	CN_out_sig(4066);
VN_in_sig(2263)	<=	CN_out_sig(4067);
VN_in_sig(3235)	<=	CN_out_sig(4068);
VN_in_sig(3783)	<=	CN_out_sig(4069);
VN_in_sig(4119)	<=	CN_out_sig(4070);
VN_in_sig(4803)	<=	CN_out_sig(4071);
VN_in_sig(523)	<=	CN_out_sig(4072);
VN_in_sig(1187)	<=	CN_out_sig(4073);
VN_in_sig(1927)	<=	CN_out_sig(4074);
VN_in_sig(2267)	<=	CN_out_sig(4075);
VN_in_sig(3239)	<=	CN_out_sig(4076);
VN_in_sig(3787)	<=	CN_out_sig(4077);
VN_in_sig(4123)	<=	CN_out_sig(4078);
VN_in_sig(4807)	<=	CN_out_sig(4079);
VN_in_sig(527)	<=	CN_out_sig(4080);
VN_in_sig(1191)	<=	CN_out_sig(4081);
VN_in_sig(1931)	<=	CN_out_sig(4082);
VN_in_sig(2271)	<=	CN_out_sig(4083);
VN_in_sig(3027)	<=	CN_out_sig(4084);
VN_in_sig(3791)	<=	CN_out_sig(4085);
VN_in_sig(4127)	<=	CN_out_sig(4086);
VN_in_sig(4811)	<=	CN_out_sig(4087);
VN_in_sig(531)	<=	CN_out_sig(4088);
VN_in_sig(1195)	<=	CN_out_sig(4089);
VN_in_sig(1935)	<=	CN_out_sig(4090);
VN_in_sig(2275)	<=	CN_out_sig(4091);
VN_in_sig(3031)	<=	CN_out_sig(4092);
VN_in_sig(3795)	<=	CN_out_sig(4093);
VN_in_sig(4131)	<=	CN_out_sig(4094);
VN_in_sig(4815)	<=	CN_out_sig(4095);
VN_in_sig(535)	<=	CN_out_sig(4096);
VN_in_sig(1199)	<=	CN_out_sig(4097);
VN_in_sig(1939)	<=	CN_out_sig(4098);
VN_in_sig(2279)	<=	CN_out_sig(4099);
VN_in_sig(3035)	<=	CN_out_sig(4100);
VN_in_sig(3799)	<=	CN_out_sig(4101);
VN_in_sig(4135)	<=	CN_out_sig(4102);
VN_in_sig(4819)	<=	CN_out_sig(4103);
VN_in_sig(539)	<=	CN_out_sig(4104);
VN_in_sig(1203)	<=	CN_out_sig(4105);
VN_in_sig(1943)	<=	CN_out_sig(4106);
VN_in_sig(2283)	<=	CN_out_sig(4107);
VN_in_sig(3039)	<=	CN_out_sig(4108);
VN_in_sig(3803)	<=	CN_out_sig(4109);
VN_in_sig(4139)	<=	CN_out_sig(4110);
VN_in_sig(4823)	<=	CN_out_sig(4111);
VN_in_sig(543)	<=	CN_out_sig(4112);
VN_in_sig(1207)	<=	CN_out_sig(4113);
VN_in_sig(1731)	<=	CN_out_sig(4114);
VN_in_sig(2287)	<=	CN_out_sig(4115);
VN_in_sig(3043)	<=	CN_out_sig(4116);
VN_in_sig(3807)	<=	CN_out_sig(4117);
VN_in_sig(4143)	<=	CN_out_sig(4118);
VN_in_sig(4827)	<=	CN_out_sig(4119);
VN_in_sig(547)	<=	CN_out_sig(4120);
VN_in_sig(1211)	<=	CN_out_sig(4121);
VN_in_sig(1735)	<=	CN_out_sig(4122);
VN_in_sig(2291)	<=	CN_out_sig(4123);
VN_in_sig(3047)	<=	CN_out_sig(4124);
VN_in_sig(3811)	<=	CN_out_sig(4125);
VN_in_sig(4147)	<=	CN_out_sig(4126);
VN_in_sig(4831)	<=	CN_out_sig(4127);
VN_in_sig(551)	<=	CN_out_sig(4128);
VN_in_sig(1215)	<=	CN_out_sig(4129);
VN_in_sig(1739)	<=	CN_out_sig(4130);
VN_in_sig(2295)	<=	CN_out_sig(4131);
VN_in_sig(3051)	<=	CN_out_sig(4132);
VN_in_sig(3815)	<=	CN_out_sig(4133);
VN_in_sig(4151)	<=	CN_out_sig(4134);
VN_in_sig(4835)	<=	CN_out_sig(4135);
VN_in_sig(555)	<=	CN_out_sig(4136);
VN_in_sig(1219)	<=	CN_out_sig(4137);
VN_in_sig(1743)	<=	CN_out_sig(4138);
VN_in_sig(2299)	<=	CN_out_sig(4139);
VN_in_sig(3055)	<=	CN_out_sig(4140);
VN_in_sig(3819)	<=	CN_out_sig(4141);
VN_in_sig(4155)	<=	CN_out_sig(4142);
VN_in_sig(4839)	<=	CN_out_sig(4143);
VN_in_sig(559)	<=	CN_out_sig(4144);
VN_in_sig(1223)	<=	CN_out_sig(4145);
VN_in_sig(1747)	<=	CN_out_sig(4146);
VN_in_sig(2303)	<=	CN_out_sig(4147);
VN_in_sig(3059)	<=	CN_out_sig(4148);
VN_in_sig(3823)	<=	CN_out_sig(4149);
VN_in_sig(4159)	<=	CN_out_sig(4150);
VN_in_sig(4843)	<=	CN_out_sig(4151);
VN_in_sig(563)	<=	CN_out_sig(4152);
VN_in_sig(1227)	<=	CN_out_sig(4153);
VN_in_sig(1751)	<=	CN_out_sig(4154);
VN_in_sig(2307)	<=	CN_out_sig(4155);
VN_in_sig(3063)	<=	CN_out_sig(4156);
VN_in_sig(3827)	<=	CN_out_sig(4157);
VN_in_sig(4163)	<=	CN_out_sig(4158);
VN_in_sig(4847)	<=	CN_out_sig(4159);
VN_in_sig(567)	<=	CN_out_sig(4160);
VN_in_sig(1231)	<=	CN_out_sig(4161);
VN_in_sig(1755)	<=	CN_out_sig(4162);
VN_in_sig(2311)	<=	CN_out_sig(4163);
VN_in_sig(3067)	<=	CN_out_sig(4164);
VN_in_sig(3831)	<=	CN_out_sig(4165);
VN_in_sig(4167)	<=	CN_out_sig(4166);
VN_in_sig(4851)	<=	CN_out_sig(4167);
VN_in_sig(571)	<=	CN_out_sig(4168);
VN_in_sig(1235)	<=	CN_out_sig(4169);
VN_in_sig(1759)	<=	CN_out_sig(4170);
VN_in_sig(2315)	<=	CN_out_sig(4171);
VN_in_sig(3071)	<=	CN_out_sig(4172);
VN_in_sig(3835)	<=	CN_out_sig(4173);
VN_in_sig(4171)	<=	CN_out_sig(4174);
VN_in_sig(4855)	<=	CN_out_sig(4175);
VN_in_sig(575)	<=	CN_out_sig(4176);
VN_in_sig(1239)	<=	CN_out_sig(4177);
VN_in_sig(1763)	<=	CN_out_sig(4178);
VN_in_sig(2319)	<=	CN_out_sig(4179);
VN_in_sig(3075)	<=	CN_out_sig(4180);
VN_in_sig(3839)	<=	CN_out_sig(4181);
VN_in_sig(4175)	<=	CN_out_sig(4182);
VN_in_sig(4859)	<=	CN_out_sig(4183);
VN_in_sig(579)	<=	CN_out_sig(4184);
VN_in_sig(1243)	<=	CN_out_sig(4185);
VN_in_sig(1767)	<=	CN_out_sig(4186);
VN_in_sig(2323)	<=	CN_out_sig(4187);
VN_in_sig(3079)	<=	CN_out_sig(4188);
VN_in_sig(3843)	<=	CN_out_sig(4189);
VN_in_sig(4179)	<=	CN_out_sig(4190);
VN_in_sig(4863)	<=	CN_out_sig(4191);
VN_in_sig(583)	<=	CN_out_sig(4192);
VN_in_sig(1247)	<=	CN_out_sig(4193);
VN_in_sig(1771)	<=	CN_out_sig(4194);
VN_in_sig(2327)	<=	CN_out_sig(4195);
VN_in_sig(3083)	<=	CN_out_sig(4196);
VN_in_sig(3847)	<=	CN_out_sig(4197);
VN_in_sig(4183)	<=	CN_out_sig(4198);
VN_in_sig(4867)	<=	CN_out_sig(4199);
VN_in_sig(587)	<=	CN_out_sig(4200);
VN_in_sig(1251)	<=	CN_out_sig(4201);
VN_in_sig(1775)	<=	CN_out_sig(4202);
VN_in_sig(2331)	<=	CN_out_sig(4203);
VN_in_sig(3087)	<=	CN_out_sig(4204);
VN_in_sig(3851)	<=	CN_out_sig(4205);
VN_in_sig(4187)	<=	CN_out_sig(4206);
VN_in_sig(4871)	<=	CN_out_sig(4207);
VN_in_sig(591)	<=	CN_out_sig(4208);
VN_in_sig(1255)	<=	CN_out_sig(4209);
VN_in_sig(1779)	<=	CN_out_sig(4210);
VN_in_sig(2335)	<=	CN_out_sig(4211);
VN_in_sig(3091)	<=	CN_out_sig(4212);
VN_in_sig(3855)	<=	CN_out_sig(4213);
VN_in_sig(4191)	<=	CN_out_sig(4214);
VN_in_sig(4875)	<=	CN_out_sig(4215);
VN_in_sig(595)	<=	CN_out_sig(4216);
VN_in_sig(1259)	<=	CN_out_sig(4217);
VN_in_sig(1783)	<=	CN_out_sig(4218);
VN_in_sig(2339)	<=	CN_out_sig(4219);
VN_in_sig(3095)	<=	CN_out_sig(4220);
VN_in_sig(3859)	<=	CN_out_sig(4221);
VN_in_sig(4195)	<=	CN_out_sig(4222);
VN_in_sig(4879)	<=	CN_out_sig(4223);
VN_in_sig(599)	<=	CN_out_sig(4224);
VN_in_sig(1263)	<=	CN_out_sig(4225);
VN_in_sig(1787)	<=	CN_out_sig(4226);
VN_in_sig(2343)	<=	CN_out_sig(4227);
VN_in_sig(3099)	<=	CN_out_sig(4228);
VN_in_sig(3863)	<=	CN_out_sig(4229);
VN_in_sig(4199)	<=	CN_out_sig(4230);
VN_in_sig(4883)	<=	CN_out_sig(4231);
VN_in_sig(603)	<=	CN_out_sig(4232);
VN_in_sig(1267)	<=	CN_out_sig(4233);
VN_in_sig(1791)	<=	CN_out_sig(4234);
VN_in_sig(2347)	<=	CN_out_sig(4235);
VN_in_sig(3103)	<=	CN_out_sig(4236);
VN_in_sig(3867)	<=	CN_out_sig(4237);
VN_in_sig(4203)	<=	CN_out_sig(4238);
VN_in_sig(4887)	<=	CN_out_sig(4239);
VN_in_sig(607)	<=	CN_out_sig(4240);
VN_in_sig(1271)	<=	CN_out_sig(4241);
VN_in_sig(1795)	<=	CN_out_sig(4242);
VN_in_sig(2351)	<=	CN_out_sig(4243);
VN_in_sig(3107)	<=	CN_out_sig(4244);
VN_in_sig(3871)	<=	CN_out_sig(4245);
VN_in_sig(4207)	<=	CN_out_sig(4246);
VN_in_sig(4891)	<=	CN_out_sig(4247);
VN_in_sig(611)	<=	CN_out_sig(4248);
VN_in_sig(1275)	<=	CN_out_sig(4249);
VN_in_sig(1799)	<=	CN_out_sig(4250);
VN_in_sig(2355)	<=	CN_out_sig(4251);
VN_in_sig(3111)	<=	CN_out_sig(4252);
VN_in_sig(3875)	<=	CN_out_sig(4253);
VN_in_sig(4211)	<=	CN_out_sig(4254);
VN_in_sig(4895)	<=	CN_out_sig(4255);
VN_in_sig(615)	<=	CN_out_sig(4256);
VN_in_sig(1279)	<=	CN_out_sig(4257);
VN_in_sig(1803)	<=	CN_out_sig(4258);
VN_in_sig(2359)	<=	CN_out_sig(4259);
VN_in_sig(3115)	<=	CN_out_sig(4260);
VN_in_sig(3879)	<=	CN_out_sig(4261);
VN_in_sig(4215)	<=	CN_out_sig(4262);
VN_in_sig(4899)	<=	CN_out_sig(4263);
VN_in_sig(619)	<=	CN_out_sig(4264);
VN_in_sig(1283)	<=	CN_out_sig(4265);
VN_in_sig(1807)	<=	CN_out_sig(4266);
VN_in_sig(2363)	<=	CN_out_sig(4267);
VN_in_sig(3119)	<=	CN_out_sig(4268);
VN_in_sig(3883)	<=	CN_out_sig(4269);
VN_in_sig(4219)	<=	CN_out_sig(4270);
VN_in_sig(4903)	<=	CN_out_sig(4271);
VN_in_sig(623)	<=	CN_out_sig(4272);
VN_in_sig(1287)	<=	CN_out_sig(4273);
VN_in_sig(1811)	<=	CN_out_sig(4274);
VN_in_sig(2367)	<=	CN_out_sig(4275);
VN_in_sig(3123)	<=	CN_out_sig(4276);
VN_in_sig(3887)	<=	CN_out_sig(4277);
VN_in_sig(4223)	<=	CN_out_sig(4278);
VN_in_sig(4907)	<=	CN_out_sig(4279);
VN_in_sig(627)	<=	CN_out_sig(4280);
VN_in_sig(1291)	<=	CN_out_sig(4281);
VN_in_sig(1815)	<=	CN_out_sig(4282);
VN_in_sig(2371)	<=	CN_out_sig(4283);
VN_in_sig(3127)	<=	CN_out_sig(4284);
VN_in_sig(3675)	<=	CN_out_sig(4285);
VN_in_sig(4227)	<=	CN_out_sig(4286);
VN_in_sig(4911)	<=	CN_out_sig(4287);
VN_in_sig(631)	<=	CN_out_sig(4288);
VN_in_sig(1295)	<=	CN_out_sig(4289);
VN_in_sig(1819)	<=	CN_out_sig(4290);
VN_in_sig(2375)	<=	CN_out_sig(4291);
VN_in_sig(3131)	<=	CN_out_sig(4292);
VN_in_sig(3679)	<=	CN_out_sig(4293);
VN_in_sig(4231)	<=	CN_out_sig(4294);
VN_in_sig(4915)	<=	CN_out_sig(4295);
VN_in_sig(635)	<=	CN_out_sig(4296);
VN_in_sig(1083)	<=	CN_out_sig(4297);
VN_in_sig(1823)	<=	CN_out_sig(4298);
VN_in_sig(2163)	<=	CN_out_sig(4299);
VN_in_sig(3135)	<=	CN_out_sig(4300);
VN_in_sig(3683)	<=	CN_out_sig(4301);
VN_in_sig(4235)	<=	CN_out_sig(4302);
VN_in_sig(4919)	<=	CN_out_sig(4303);
VN_in_sig(639)	<=	CN_out_sig(4304);
VN_in_sig(1087)	<=	CN_out_sig(4305);
VN_in_sig(1827)	<=	CN_out_sig(4306);
VN_in_sig(2167)	<=	CN_out_sig(4307);
VN_in_sig(3139)	<=	CN_out_sig(4308);
VN_in_sig(3687)	<=	CN_out_sig(4309);
VN_in_sig(4239)	<=	CN_out_sig(4310);
VN_in_sig(4923)	<=	CN_out_sig(4311);
VN_in_sig(643)	<=	CN_out_sig(4312);
VN_in_sig(1091)	<=	CN_out_sig(4313);
VN_in_sig(1831)	<=	CN_out_sig(4314);
VN_in_sig(2171)	<=	CN_out_sig(4315);
VN_in_sig(3143)	<=	CN_out_sig(4316);
VN_in_sig(3691)	<=	CN_out_sig(4317);
VN_in_sig(4243)	<=	CN_out_sig(4318);
VN_in_sig(4927)	<=	CN_out_sig(4319);
VN_in_sig(235)	<=	CN_out_sig(4320);
VN_in_sig(883)	<=	CN_out_sig(4321);
VN_in_sig(1535)	<=	CN_out_sig(4322);
VN_in_sig(2431)	<=	CN_out_sig(4323);
VN_in_sig(2763)	<=	CN_out_sig(4324);
VN_in_sig(3443)	<=	CN_out_sig(4325);
VN_in_sig(4467)	<=	CN_out_sig(4326);
VN_in_sig(4691)	<=	CN_out_sig(4327);
VN_in_sig(239)	<=	CN_out_sig(4328);
VN_in_sig(887)	<=	CN_out_sig(4329);
VN_in_sig(1539)	<=	CN_out_sig(4330);
VN_in_sig(2435)	<=	CN_out_sig(4331);
VN_in_sig(2767)	<=	CN_out_sig(4332);
VN_in_sig(3447)	<=	CN_out_sig(4333);
VN_in_sig(4471)	<=	CN_out_sig(4334);
VN_in_sig(4695)	<=	CN_out_sig(4335);
VN_in_sig(243)	<=	CN_out_sig(4336);
VN_in_sig(891)	<=	CN_out_sig(4337);
VN_in_sig(1543)	<=	CN_out_sig(4338);
VN_in_sig(2439)	<=	CN_out_sig(4339);
VN_in_sig(2771)	<=	CN_out_sig(4340);
VN_in_sig(3451)	<=	CN_out_sig(4341);
VN_in_sig(4475)	<=	CN_out_sig(4342);
VN_in_sig(4699)	<=	CN_out_sig(4343);
VN_in_sig(247)	<=	CN_out_sig(4344);
VN_in_sig(895)	<=	CN_out_sig(4345);
VN_in_sig(1547)	<=	CN_out_sig(4346);
VN_in_sig(2443)	<=	CN_out_sig(4347);
VN_in_sig(2775)	<=	CN_out_sig(4348);
VN_in_sig(3455)	<=	CN_out_sig(4349);
VN_in_sig(4479)	<=	CN_out_sig(4350);
VN_in_sig(4703)	<=	CN_out_sig(4351);
VN_in_sig(251)	<=	CN_out_sig(4352);
VN_in_sig(899)	<=	CN_out_sig(4353);
VN_in_sig(1551)	<=	CN_out_sig(4354);
VN_in_sig(2447)	<=	CN_out_sig(4355);
VN_in_sig(2779)	<=	CN_out_sig(4356);
VN_in_sig(3243)	<=	CN_out_sig(4357);
VN_in_sig(4483)	<=	CN_out_sig(4358);
VN_in_sig(4707)	<=	CN_out_sig(4359);
VN_in_sig(255)	<=	CN_out_sig(4360);
VN_in_sig(903)	<=	CN_out_sig(4361);
VN_in_sig(1555)	<=	CN_out_sig(4362);
VN_in_sig(2451)	<=	CN_out_sig(4363);
VN_in_sig(2783)	<=	CN_out_sig(4364);
VN_in_sig(3247)	<=	CN_out_sig(4365);
VN_in_sig(4487)	<=	CN_out_sig(4366);
VN_in_sig(4711)	<=	CN_out_sig(4367);
VN_in_sig(259)	<=	CN_out_sig(4368);
VN_in_sig(907)	<=	CN_out_sig(4369);
VN_in_sig(1559)	<=	CN_out_sig(4370);
VN_in_sig(2455)	<=	CN_out_sig(4371);
VN_in_sig(2787)	<=	CN_out_sig(4372);
VN_in_sig(3251)	<=	CN_out_sig(4373);
VN_in_sig(4491)	<=	CN_out_sig(4374);
VN_in_sig(4715)	<=	CN_out_sig(4375);
VN_in_sig(263)	<=	CN_out_sig(4376);
VN_in_sig(911)	<=	CN_out_sig(4377);
VN_in_sig(1563)	<=	CN_out_sig(4378);
VN_in_sig(2459)	<=	CN_out_sig(4379);
VN_in_sig(2791)	<=	CN_out_sig(4380);
VN_in_sig(3255)	<=	CN_out_sig(4381);
VN_in_sig(4495)	<=	CN_out_sig(4382);
VN_in_sig(4719)	<=	CN_out_sig(4383);
VN_in_sig(267)	<=	CN_out_sig(4384);
VN_in_sig(915)	<=	CN_out_sig(4385);
VN_in_sig(1567)	<=	CN_out_sig(4386);
VN_in_sig(2463)	<=	CN_out_sig(4387);
VN_in_sig(2795)	<=	CN_out_sig(4388);
VN_in_sig(3259)	<=	CN_out_sig(4389);
VN_in_sig(4499)	<=	CN_out_sig(4390);
VN_in_sig(4723)	<=	CN_out_sig(4391);
VN_in_sig(271)	<=	CN_out_sig(4392);
VN_in_sig(919)	<=	CN_out_sig(4393);
VN_in_sig(1571)	<=	CN_out_sig(4394);
VN_in_sig(2467)	<=	CN_out_sig(4395);
VN_in_sig(2799)	<=	CN_out_sig(4396);
VN_in_sig(3263)	<=	CN_out_sig(4397);
VN_in_sig(4503)	<=	CN_out_sig(4398);
VN_in_sig(4727)	<=	CN_out_sig(4399);
VN_in_sig(275)	<=	CN_out_sig(4400);
VN_in_sig(923)	<=	CN_out_sig(4401);
VN_in_sig(1575)	<=	CN_out_sig(4402);
VN_in_sig(2471)	<=	CN_out_sig(4403);
VN_in_sig(2803)	<=	CN_out_sig(4404);
VN_in_sig(3267)	<=	CN_out_sig(4405);
VN_in_sig(4507)	<=	CN_out_sig(4406);
VN_in_sig(4731)	<=	CN_out_sig(4407);
VN_in_sig(279)	<=	CN_out_sig(4408);
VN_in_sig(927)	<=	CN_out_sig(4409);
VN_in_sig(1579)	<=	CN_out_sig(4410);
VN_in_sig(2475)	<=	CN_out_sig(4411);
VN_in_sig(2807)	<=	CN_out_sig(4412);
VN_in_sig(3271)	<=	CN_out_sig(4413);
VN_in_sig(4511)	<=	CN_out_sig(4414);
VN_in_sig(4735)	<=	CN_out_sig(4415);
VN_in_sig(283)	<=	CN_out_sig(4416);
VN_in_sig(931)	<=	CN_out_sig(4417);
VN_in_sig(1583)	<=	CN_out_sig(4418);
VN_in_sig(2479)	<=	CN_out_sig(4419);
VN_in_sig(2595)	<=	CN_out_sig(4420);
VN_in_sig(3275)	<=	CN_out_sig(4421);
VN_in_sig(4515)	<=	CN_out_sig(4422);
VN_in_sig(4739)	<=	CN_out_sig(4423);
VN_in_sig(287)	<=	CN_out_sig(4424);
VN_in_sig(935)	<=	CN_out_sig(4425);
VN_in_sig(1587)	<=	CN_out_sig(4426);
VN_in_sig(2483)	<=	CN_out_sig(4427);
VN_in_sig(2599)	<=	CN_out_sig(4428);
VN_in_sig(3279)	<=	CN_out_sig(4429);
VN_in_sig(4519)	<=	CN_out_sig(4430);
VN_in_sig(4743)	<=	CN_out_sig(4431);
VN_in_sig(291)	<=	CN_out_sig(4432);
VN_in_sig(939)	<=	CN_out_sig(4433);
VN_in_sig(1591)	<=	CN_out_sig(4434);
VN_in_sig(2487)	<=	CN_out_sig(4435);
VN_in_sig(2603)	<=	CN_out_sig(4436);
VN_in_sig(3283)	<=	CN_out_sig(4437);
VN_in_sig(4523)	<=	CN_out_sig(4438);
VN_in_sig(4747)	<=	CN_out_sig(4439);
VN_in_sig(295)	<=	CN_out_sig(4440);
VN_in_sig(943)	<=	CN_out_sig(4441);
VN_in_sig(1595)	<=	CN_out_sig(4442);
VN_in_sig(2491)	<=	CN_out_sig(4443);
VN_in_sig(2607)	<=	CN_out_sig(4444);
VN_in_sig(3287)	<=	CN_out_sig(4445);
VN_in_sig(4527)	<=	CN_out_sig(4446);
VN_in_sig(4751)	<=	CN_out_sig(4447);
VN_in_sig(299)	<=	CN_out_sig(4448);
VN_in_sig(947)	<=	CN_out_sig(4449);
VN_in_sig(1599)	<=	CN_out_sig(4450);
VN_in_sig(2495)	<=	CN_out_sig(4451);
VN_in_sig(2611)	<=	CN_out_sig(4452);
VN_in_sig(3291)	<=	CN_out_sig(4453);
VN_in_sig(4531)	<=	CN_out_sig(4454);
VN_in_sig(4539)	<=	CN_out_sig(4455);
VN_in_sig(303)	<=	CN_out_sig(4456);
VN_in_sig(951)	<=	CN_out_sig(4457);
VN_in_sig(1603)	<=	CN_out_sig(4458);
VN_in_sig(2499)	<=	CN_out_sig(4459);
VN_in_sig(2615)	<=	CN_out_sig(4460);
VN_in_sig(3295)	<=	CN_out_sig(4461);
VN_in_sig(4535)	<=	CN_out_sig(4462);
VN_in_sig(4543)	<=	CN_out_sig(4463);
VN_in_sig(307)	<=	CN_out_sig(4464);
VN_in_sig(955)	<=	CN_out_sig(4465);
VN_in_sig(1607)	<=	CN_out_sig(4466);
VN_in_sig(2503)	<=	CN_out_sig(4467);
VN_in_sig(2619)	<=	CN_out_sig(4468);
VN_in_sig(3299)	<=	CN_out_sig(4469);
VN_in_sig(4323)	<=	CN_out_sig(4470);
VN_in_sig(4547)	<=	CN_out_sig(4471);
VN_in_sig(311)	<=	CN_out_sig(4472);
VN_in_sig(959)	<=	CN_out_sig(4473);
VN_in_sig(1611)	<=	CN_out_sig(4474);
VN_in_sig(2507)	<=	CN_out_sig(4475);
VN_in_sig(2623)	<=	CN_out_sig(4476);
VN_in_sig(3303)	<=	CN_out_sig(4477);
VN_in_sig(4327)	<=	CN_out_sig(4478);
VN_in_sig(4551)	<=	CN_out_sig(4479);
VN_in_sig(315)	<=	CN_out_sig(4480);
VN_in_sig(963)	<=	CN_out_sig(4481);
VN_in_sig(1615)	<=	CN_out_sig(4482);
VN_in_sig(2511)	<=	CN_out_sig(4483);
VN_in_sig(2627)	<=	CN_out_sig(4484);
VN_in_sig(3307)	<=	CN_out_sig(4485);
VN_in_sig(4331)	<=	CN_out_sig(4486);
VN_in_sig(4555)	<=	CN_out_sig(4487);
VN_in_sig(319)	<=	CN_out_sig(4488);
VN_in_sig(967)	<=	CN_out_sig(4489);
VN_in_sig(1619)	<=	CN_out_sig(4490);
VN_in_sig(2515)	<=	CN_out_sig(4491);
VN_in_sig(2631)	<=	CN_out_sig(4492);
VN_in_sig(3311)	<=	CN_out_sig(4493);
VN_in_sig(4335)	<=	CN_out_sig(4494);
VN_in_sig(4559)	<=	CN_out_sig(4495);
VN_in_sig(323)	<=	CN_out_sig(4496);
VN_in_sig(971)	<=	CN_out_sig(4497);
VN_in_sig(1623)	<=	CN_out_sig(4498);
VN_in_sig(2519)	<=	CN_out_sig(4499);
VN_in_sig(2635)	<=	CN_out_sig(4500);
VN_in_sig(3315)	<=	CN_out_sig(4501);
VN_in_sig(4339)	<=	CN_out_sig(4502);
VN_in_sig(4563)	<=	CN_out_sig(4503);
VN_in_sig(327)	<=	CN_out_sig(4504);
VN_in_sig(975)	<=	CN_out_sig(4505);
VN_in_sig(1627)	<=	CN_out_sig(4506);
VN_in_sig(2523)	<=	CN_out_sig(4507);
VN_in_sig(2639)	<=	CN_out_sig(4508);
VN_in_sig(3319)	<=	CN_out_sig(4509);
VN_in_sig(4343)	<=	CN_out_sig(4510);
VN_in_sig(4567)	<=	CN_out_sig(4511);
VN_in_sig(331)	<=	CN_out_sig(4512);
VN_in_sig(979)	<=	CN_out_sig(4513);
VN_in_sig(1631)	<=	CN_out_sig(4514);
VN_in_sig(2527)	<=	CN_out_sig(4515);
VN_in_sig(2643)	<=	CN_out_sig(4516);
VN_in_sig(3323)	<=	CN_out_sig(4517);
VN_in_sig(4347)	<=	CN_out_sig(4518);
VN_in_sig(4571)	<=	CN_out_sig(4519);
VN_in_sig(335)	<=	CN_out_sig(4520);
VN_in_sig(983)	<=	CN_out_sig(4521);
VN_in_sig(1635)	<=	CN_out_sig(4522);
VN_in_sig(2531)	<=	CN_out_sig(4523);
VN_in_sig(2647)	<=	CN_out_sig(4524);
VN_in_sig(3327)	<=	CN_out_sig(4525);
VN_in_sig(4351)	<=	CN_out_sig(4526);
VN_in_sig(4575)	<=	CN_out_sig(4527);
VN_in_sig(339)	<=	CN_out_sig(4528);
VN_in_sig(987)	<=	CN_out_sig(4529);
VN_in_sig(1639)	<=	CN_out_sig(4530);
VN_in_sig(2535)	<=	CN_out_sig(4531);
VN_in_sig(2651)	<=	CN_out_sig(4532);
VN_in_sig(3331)	<=	CN_out_sig(4533);
VN_in_sig(4355)	<=	CN_out_sig(4534);
VN_in_sig(4579)	<=	CN_out_sig(4535);
VN_in_sig(343)	<=	CN_out_sig(4536);
VN_in_sig(991)	<=	CN_out_sig(4537);
VN_in_sig(1643)	<=	CN_out_sig(4538);
VN_in_sig(2539)	<=	CN_out_sig(4539);
VN_in_sig(2655)	<=	CN_out_sig(4540);
VN_in_sig(3335)	<=	CN_out_sig(4541);
VN_in_sig(4359)	<=	CN_out_sig(4542);
VN_in_sig(4583)	<=	CN_out_sig(4543);
VN_in_sig(347)	<=	CN_out_sig(4544);
VN_in_sig(995)	<=	CN_out_sig(4545);
VN_in_sig(1647)	<=	CN_out_sig(4546);
VN_in_sig(2543)	<=	CN_out_sig(4547);
VN_in_sig(2659)	<=	CN_out_sig(4548);
VN_in_sig(3339)	<=	CN_out_sig(4549);
VN_in_sig(4363)	<=	CN_out_sig(4550);
VN_in_sig(4587)	<=	CN_out_sig(4551);
VN_in_sig(351)	<=	CN_out_sig(4552);
VN_in_sig(999)	<=	CN_out_sig(4553);
VN_in_sig(1651)	<=	CN_out_sig(4554);
VN_in_sig(2547)	<=	CN_out_sig(4555);
VN_in_sig(2663)	<=	CN_out_sig(4556);
VN_in_sig(3343)	<=	CN_out_sig(4557);
VN_in_sig(4367)	<=	CN_out_sig(4558);
VN_in_sig(4591)	<=	CN_out_sig(4559);
VN_in_sig(355)	<=	CN_out_sig(4560);
VN_in_sig(1003)	<=	CN_out_sig(4561);
VN_in_sig(1655)	<=	CN_out_sig(4562);
VN_in_sig(2551)	<=	CN_out_sig(4563);
VN_in_sig(2667)	<=	CN_out_sig(4564);
VN_in_sig(3347)	<=	CN_out_sig(4565);
VN_in_sig(4371)	<=	CN_out_sig(4566);
VN_in_sig(4595)	<=	CN_out_sig(4567);
VN_in_sig(359)	<=	CN_out_sig(4568);
VN_in_sig(1007)	<=	CN_out_sig(4569);
VN_in_sig(1659)	<=	CN_out_sig(4570);
VN_in_sig(2555)	<=	CN_out_sig(4571);
VN_in_sig(2671)	<=	CN_out_sig(4572);
VN_in_sig(3351)	<=	CN_out_sig(4573);
VN_in_sig(4375)	<=	CN_out_sig(4574);
VN_in_sig(4599)	<=	CN_out_sig(4575);
VN_in_sig(363)	<=	CN_out_sig(4576);
VN_in_sig(1011)	<=	CN_out_sig(4577);
VN_in_sig(1663)	<=	CN_out_sig(4578);
VN_in_sig(2559)	<=	CN_out_sig(4579);
VN_in_sig(2675)	<=	CN_out_sig(4580);
VN_in_sig(3355)	<=	CN_out_sig(4581);
VN_in_sig(4379)	<=	CN_out_sig(4582);
VN_in_sig(4603)	<=	CN_out_sig(4583);
VN_in_sig(367)	<=	CN_out_sig(4584);
VN_in_sig(1015)	<=	CN_out_sig(4585);
VN_in_sig(1667)	<=	CN_out_sig(4586);
VN_in_sig(2563)	<=	CN_out_sig(4587);
VN_in_sig(2679)	<=	CN_out_sig(4588);
VN_in_sig(3359)	<=	CN_out_sig(4589);
VN_in_sig(4383)	<=	CN_out_sig(4590);
VN_in_sig(4607)	<=	CN_out_sig(4591);
VN_in_sig(371)	<=	CN_out_sig(4592);
VN_in_sig(1019)	<=	CN_out_sig(4593);
VN_in_sig(1671)	<=	CN_out_sig(4594);
VN_in_sig(2567)	<=	CN_out_sig(4595);
VN_in_sig(2683)	<=	CN_out_sig(4596);
VN_in_sig(3363)	<=	CN_out_sig(4597);
VN_in_sig(4387)	<=	CN_out_sig(4598);
VN_in_sig(4611)	<=	CN_out_sig(4599);
VN_in_sig(375)	<=	CN_out_sig(4600);
VN_in_sig(1023)	<=	CN_out_sig(4601);
VN_in_sig(1675)	<=	CN_out_sig(4602);
VN_in_sig(2571)	<=	CN_out_sig(4603);
VN_in_sig(2687)	<=	CN_out_sig(4604);
VN_in_sig(3367)	<=	CN_out_sig(4605);
VN_in_sig(4391)	<=	CN_out_sig(4606);
VN_in_sig(4615)	<=	CN_out_sig(4607);
VN_in_sig(379)	<=	CN_out_sig(4608);
VN_in_sig(1027)	<=	CN_out_sig(4609);
VN_in_sig(1679)	<=	CN_out_sig(4610);
VN_in_sig(2575)	<=	CN_out_sig(4611);
VN_in_sig(2691)	<=	CN_out_sig(4612);
VN_in_sig(3371)	<=	CN_out_sig(4613);
VN_in_sig(4395)	<=	CN_out_sig(4614);
VN_in_sig(4619)	<=	CN_out_sig(4615);
VN_in_sig(383)	<=	CN_out_sig(4616);
VN_in_sig(1031)	<=	CN_out_sig(4617);
VN_in_sig(1683)	<=	CN_out_sig(4618);
VN_in_sig(2579)	<=	CN_out_sig(4619);
VN_in_sig(2695)	<=	CN_out_sig(4620);
VN_in_sig(3375)	<=	CN_out_sig(4621);
VN_in_sig(4399)	<=	CN_out_sig(4622);
VN_in_sig(4623)	<=	CN_out_sig(4623);
VN_in_sig(387)	<=	CN_out_sig(4624);
VN_in_sig(1035)	<=	CN_out_sig(4625);
VN_in_sig(1687)	<=	CN_out_sig(4626);
VN_in_sig(2583)	<=	CN_out_sig(4627);
VN_in_sig(2699)	<=	CN_out_sig(4628);
VN_in_sig(3379)	<=	CN_out_sig(4629);
VN_in_sig(4403)	<=	CN_out_sig(4630);
VN_in_sig(4627)	<=	CN_out_sig(4631);
VN_in_sig(391)	<=	CN_out_sig(4632);
VN_in_sig(1039)	<=	CN_out_sig(4633);
VN_in_sig(1691)	<=	CN_out_sig(4634);
VN_in_sig(2587)	<=	CN_out_sig(4635);
VN_in_sig(2703)	<=	CN_out_sig(4636);
VN_in_sig(3383)	<=	CN_out_sig(4637);
VN_in_sig(4407)	<=	CN_out_sig(4638);
VN_in_sig(4631)	<=	CN_out_sig(4639);
VN_in_sig(395)	<=	CN_out_sig(4640);
VN_in_sig(1043)	<=	CN_out_sig(4641);
VN_in_sig(1695)	<=	CN_out_sig(4642);
VN_in_sig(2591)	<=	CN_out_sig(4643);
VN_in_sig(2707)	<=	CN_out_sig(4644);
VN_in_sig(3387)	<=	CN_out_sig(4645);
VN_in_sig(4411)	<=	CN_out_sig(4646);
VN_in_sig(4635)	<=	CN_out_sig(4647);
VN_in_sig(399)	<=	CN_out_sig(4648);
VN_in_sig(1047)	<=	CN_out_sig(4649);
VN_in_sig(1699)	<=	CN_out_sig(4650);
VN_in_sig(2379)	<=	CN_out_sig(4651);
VN_in_sig(2711)	<=	CN_out_sig(4652);
VN_in_sig(3391)	<=	CN_out_sig(4653);
VN_in_sig(4415)	<=	CN_out_sig(4654);
VN_in_sig(4639)	<=	CN_out_sig(4655);
VN_in_sig(403)	<=	CN_out_sig(4656);
VN_in_sig(1051)	<=	CN_out_sig(4657);
VN_in_sig(1703)	<=	CN_out_sig(4658);
VN_in_sig(2383)	<=	CN_out_sig(4659);
VN_in_sig(2715)	<=	CN_out_sig(4660);
VN_in_sig(3395)	<=	CN_out_sig(4661);
VN_in_sig(4419)	<=	CN_out_sig(4662);
VN_in_sig(4643)	<=	CN_out_sig(4663);
VN_in_sig(407)	<=	CN_out_sig(4664);
VN_in_sig(1055)	<=	CN_out_sig(4665);
VN_in_sig(1707)	<=	CN_out_sig(4666);
VN_in_sig(2387)	<=	CN_out_sig(4667);
VN_in_sig(2719)	<=	CN_out_sig(4668);
VN_in_sig(3399)	<=	CN_out_sig(4669);
VN_in_sig(4423)	<=	CN_out_sig(4670);
VN_in_sig(4647)	<=	CN_out_sig(4671);
VN_in_sig(411)	<=	CN_out_sig(4672);
VN_in_sig(1059)	<=	CN_out_sig(4673);
VN_in_sig(1711)	<=	CN_out_sig(4674);
VN_in_sig(2391)	<=	CN_out_sig(4675);
VN_in_sig(2723)	<=	CN_out_sig(4676);
VN_in_sig(3403)	<=	CN_out_sig(4677);
VN_in_sig(4427)	<=	CN_out_sig(4678);
VN_in_sig(4651)	<=	CN_out_sig(4679);
VN_in_sig(415)	<=	CN_out_sig(4680);
VN_in_sig(1063)	<=	CN_out_sig(4681);
VN_in_sig(1715)	<=	CN_out_sig(4682);
VN_in_sig(2395)	<=	CN_out_sig(4683);
VN_in_sig(2727)	<=	CN_out_sig(4684);
VN_in_sig(3407)	<=	CN_out_sig(4685);
VN_in_sig(4431)	<=	CN_out_sig(4686);
VN_in_sig(4655)	<=	CN_out_sig(4687);
VN_in_sig(419)	<=	CN_out_sig(4688);
VN_in_sig(1067)	<=	CN_out_sig(4689);
VN_in_sig(1719)	<=	CN_out_sig(4690);
VN_in_sig(2399)	<=	CN_out_sig(4691);
VN_in_sig(2731)	<=	CN_out_sig(4692);
VN_in_sig(3411)	<=	CN_out_sig(4693);
VN_in_sig(4435)	<=	CN_out_sig(4694);
VN_in_sig(4659)	<=	CN_out_sig(4695);
VN_in_sig(423)	<=	CN_out_sig(4696);
VN_in_sig(1071)	<=	CN_out_sig(4697);
VN_in_sig(1723)	<=	CN_out_sig(4698);
VN_in_sig(2403)	<=	CN_out_sig(4699);
VN_in_sig(2735)	<=	CN_out_sig(4700);
VN_in_sig(3415)	<=	CN_out_sig(4701);
VN_in_sig(4439)	<=	CN_out_sig(4702);
VN_in_sig(4663)	<=	CN_out_sig(4703);
VN_in_sig(427)	<=	CN_out_sig(4704);
VN_in_sig(1075)	<=	CN_out_sig(4705);
VN_in_sig(1727)	<=	CN_out_sig(4706);
VN_in_sig(2407)	<=	CN_out_sig(4707);
VN_in_sig(2739)	<=	CN_out_sig(4708);
VN_in_sig(3419)	<=	CN_out_sig(4709);
VN_in_sig(4443)	<=	CN_out_sig(4710);
VN_in_sig(4667)	<=	CN_out_sig(4711);
VN_in_sig(431)	<=	CN_out_sig(4712);
VN_in_sig(1079)	<=	CN_out_sig(4713);
VN_in_sig(1515)	<=	CN_out_sig(4714);
VN_in_sig(2411)	<=	CN_out_sig(4715);
VN_in_sig(2743)	<=	CN_out_sig(4716);
VN_in_sig(3423)	<=	CN_out_sig(4717);
VN_in_sig(4447)	<=	CN_out_sig(4718);
VN_in_sig(4671)	<=	CN_out_sig(4719);
VN_in_sig(219)	<=	CN_out_sig(4720);
VN_in_sig(867)	<=	CN_out_sig(4721);
VN_in_sig(1519)	<=	CN_out_sig(4722);
VN_in_sig(2415)	<=	CN_out_sig(4723);
VN_in_sig(2747)	<=	CN_out_sig(4724);
VN_in_sig(3427)	<=	CN_out_sig(4725);
VN_in_sig(4451)	<=	CN_out_sig(4726);
VN_in_sig(4675)	<=	CN_out_sig(4727);
VN_in_sig(223)	<=	CN_out_sig(4728);
VN_in_sig(871)	<=	CN_out_sig(4729);
VN_in_sig(1523)	<=	CN_out_sig(4730);
VN_in_sig(2419)	<=	CN_out_sig(4731);
VN_in_sig(2751)	<=	CN_out_sig(4732);
VN_in_sig(3431)	<=	CN_out_sig(4733);
VN_in_sig(4455)	<=	CN_out_sig(4734);
VN_in_sig(4679)	<=	CN_out_sig(4735);
VN_in_sig(227)	<=	CN_out_sig(4736);
VN_in_sig(875)	<=	CN_out_sig(4737);
VN_in_sig(1527)	<=	CN_out_sig(4738);
VN_in_sig(2423)	<=	CN_out_sig(4739);
VN_in_sig(2755)	<=	CN_out_sig(4740);
VN_in_sig(3435)	<=	CN_out_sig(4741);
VN_in_sig(4459)	<=	CN_out_sig(4742);
VN_in_sig(4683)	<=	CN_out_sig(4743);
VN_in_sig(231)	<=	CN_out_sig(4744);
VN_in_sig(879)	<=	CN_out_sig(4745);
VN_in_sig(1531)	<=	CN_out_sig(4746);
VN_in_sig(2427)	<=	CN_out_sig(4747);
VN_in_sig(2759)	<=	CN_out_sig(4748);
VN_in_sig(3439)	<=	CN_out_sig(4749);
VN_in_sig(4463)	<=	CN_out_sig(4750);
VN_in_sig(4687)	<=	CN_out_sig(4751);
VN_in_sig(159)	<=	CN_out_sig(4752);
VN_in_sig(719)	<=	CN_out_sig(4753);
VN_in_sig(1443)	<=	CN_out_sig(4754);
VN_in_sig(2083)	<=	CN_out_sig(4755);
VN_in_sig(2995)	<=	CN_out_sig(4756);
VN_in_sig(3507)	<=	CN_out_sig(4757);
VN_in_sig(3923)	<=	CN_out_sig(4758);
VN_in_sig(5031)	<=	CN_out_sig(4759);
VN_in_sig(163)	<=	CN_out_sig(4760);
VN_in_sig(723)	<=	CN_out_sig(4761);
VN_in_sig(1447)	<=	CN_out_sig(4762);
VN_in_sig(2087)	<=	CN_out_sig(4763);
VN_in_sig(2999)	<=	CN_out_sig(4764);
VN_in_sig(3511)	<=	CN_out_sig(4765);
VN_in_sig(3927)	<=	CN_out_sig(4766);
VN_in_sig(5035)	<=	CN_out_sig(4767);
VN_in_sig(167)	<=	CN_out_sig(4768);
VN_in_sig(727)	<=	CN_out_sig(4769);
VN_in_sig(1451)	<=	CN_out_sig(4770);
VN_in_sig(2091)	<=	CN_out_sig(4771);
VN_in_sig(3003)	<=	CN_out_sig(4772);
VN_in_sig(3515)	<=	CN_out_sig(4773);
VN_in_sig(3931)	<=	CN_out_sig(4774);
VN_in_sig(5039)	<=	CN_out_sig(4775);
VN_in_sig(171)	<=	CN_out_sig(4776);
VN_in_sig(731)	<=	CN_out_sig(4777);
VN_in_sig(1455)	<=	CN_out_sig(4778);
VN_in_sig(2095)	<=	CN_out_sig(4779);
VN_in_sig(3007)	<=	CN_out_sig(4780);
VN_in_sig(3519)	<=	CN_out_sig(4781);
VN_in_sig(3935)	<=	CN_out_sig(4782);
VN_in_sig(5043)	<=	CN_out_sig(4783);
VN_in_sig(175)	<=	CN_out_sig(4784);
VN_in_sig(735)	<=	CN_out_sig(4785);
VN_in_sig(1459)	<=	CN_out_sig(4786);
VN_in_sig(2099)	<=	CN_out_sig(4787);
VN_in_sig(3011)	<=	CN_out_sig(4788);
VN_in_sig(3523)	<=	CN_out_sig(4789);
VN_in_sig(3939)	<=	CN_out_sig(4790);
VN_in_sig(5047)	<=	CN_out_sig(4791);
VN_in_sig(179)	<=	CN_out_sig(4792);
VN_in_sig(739)	<=	CN_out_sig(4793);
VN_in_sig(1463)	<=	CN_out_sig(4794);
VN_in_sig(2103)	<=	CN_out_sig(4795);
VN_in_sig(3015)	<=	CN_out_sig(4796);
VN_in_sig(3527)	<=	CN_out_sig(4797);
VN_in_sig(3943)	<=	CN_out_sig(4798);
VN_in_sig(5051)	<=	CN_out_sig(4799);
VN_in_sig(183)	<=	CN_out_sig(4800);
VN_in_sig(743)	<=	CN_out_sig(4801);
VN_in_sig(1467)	<=	CN_out_sig(4802);
VN_in_sig(2107)	<=	CN_out_sig(4803);
VN_in_sig(3019)	<=	CN_out_sig(4804);
VN_in_sig(3531)	<=	CN_out_sig(4805);
VN_in_sig(3947)	<=	CN_out_sig(4806);
VN_in_sig(5055)	<=	CN_out_sig(4807);
VN_in_sig(187)	<=	CN_out_sig(4808);
VN_in_sig(747)	<=	CN_out_sig(4809);
VN_in_sig(1471)	<=	CN_out_sig(4810);
VN_in_sig(2111)	<=	CN_out_sig(4811);
VN_in_sig(3023)	<=	CN_out_sig(4812);
VN_in_sig(3535)	<=	CN_out_sig(4813);
VN_in_sig(3951)	<=	CN_out_sig(4814);
VN_in_sig(5059)	<=	CN_out_sig(4815);
VN_in_sig(191)	<=	CN_out_sig(4816);
VN_in_sig(751)	<=	CN_out_sig(4817);
VN_in_sig(1475)	<=	CN_out_sig(4818);
VN_in_sig(2115)	<=	CN_out_sig(4819);
VN_in_sig(2811)	<=	CN_out_sig(4820);
VN_in_sig(3539)	<=	CN_out_sig(4821);
VN_in_sig(3955)	<=	CN_out_sig(4822);
VN_in_sig(5063)	<=	CN_out_sig(4823);
VN_in_sig(195)	<=	CN_out_sig(4824);
VN_in_sig(755)	<=	CN_out_sig(4825);
VN_in_sig(1479)	<=	CN_out_sig(4826);
VN_in_sig(2119)	<=	CN_out_sig(4827);
VN_in_sig(2815)	<=	CN_out_sig(4828);
VN_in_sig(3543)	<=	CN_out_sig(4829);
VN_in_sig(3959)	<=	CN_out_sig(4830);
VN_in_sig(5067)	<=	CN_out_sig(4831);
VN_in_sig(199)	<=	CN_out_sig(4832);
VN_in_sig(759)	<=	CN_out_sig(4833);
VN_in_sig(1483)	<=	CN_out_sig(4834);
VN_in_sig(2123)	<=	CN_out_sig(4835);
VN_in_sig(2819)	<=	CN_out_sig(4836);
VN_in_sig(3547)	<=	CN_out_sig(4837);
VN_in_sig(3963)	<=	CN_out_sig(4838);
VN_in_sig(5071)	<=	CN_out_sig(4839);
VN_in_sig(203)	<=	CN_out_sig(4840);
VN_in_sig(763)	<=	CN_out_sig(4841);
VN_in_sig(1487)	<=	CN_out_sig(4842);
VN_in_sig(2127)	<=	CN_out_sig(4843);
VN_in_sig(2823)	<=	CN_out_sig(4844);
VN_in_sig(3551)	<=	CN_out_sig(4845);
VN_in_sig(3967)	<=	CN_out_sig(4846);
VN_in_sig(5075)	<=	CN_out_sig(4847);
VN_in_sig(207)	<=	CN_out_sig(4848);
VN_in_sig(767)	<=	CN_out_sig(4849);
VN_in_sig(1491)	<=	CN_out_sig(4850);
VN_in_sig(2131)	<=	CN_out_sig(4851);
VN_in_sig(2827)	<=	CN_out_sig(4852);
VN_in_sig(3555)	<=	CN_out_sig(4853);
VN_in_sig(3971)	<=	CN_out_sig(4854);
VN_in_sig(5079)	<=	CN_out_sig(4855);
VN_in_sig(211)	<=	CN_out_sig(4856);
VN_in_sig(771)	<=	CN_out_sig(4857);
VN_in_sig(1495)	<=	CN_out_sig(4858);
VN_in_sig(2135)	<=	CN_out_sig(4859);
VN_in_sig(2831)	<=	CN_out_sig(4860);
VN_in_sig(3559)	<=	CN_out_sig(4861);
VN_in_sig(3975)	<=	CN_out_sig(4862);
VN_in_sig(5083)	<=	CN_out_sig(4863);
VN_in_sig(215)	<=	CN_out_sig(4864);
VN_in_sig(775)	<=	CN_out_sig(4865);
VN_in_sig(1499)	<=	CN_out_sig(4866);
VN_in_sig(2139)	<=	CN_out_sig(4867);
VN_in_sig(2835)	<=	CN_out_sig(4868);
VN_in_sig(3563)	<=	CN_out_sig(4869);
VN_in_sig(3979)	<=	CN_out_sig(4870);
VN_in_sig(5087)	<=	CN_out_sig(4871);
VN_in_sig(3)	<=	CN_out_sig(4872);
VN_in_sig(779)	<=	CN_out_sig(4873);
VN_in_sig(1503)	<=	CN_out_sig(4874);
VN_in_sig(2143)	<=	CN_out_sig(4875);
VN_in_sig(2839)	<=	CN_out_sig(4876);
VN_in_sig(3567)	<=	CN_out_sig(4877);
VN_in_sig(3983)	<=	CN_out_sig(4878);
VN_in_sig(5091)	<=	CN_out_sig(4879);
VN_in_sig(7)	<=	CN_out_sig(4880);
VN_in_sig(783)	<=	CN_out_sig(4881);
VN_in_sig(1507)	<=	CN_out_sig(4882);
VN_in_sig(2147)	<=	CN_out_sig(4883);
VN_in_sig(2843)	<=	CN_out_sig(4884);
VN_in_sig(3571)	<=	CN_out_sig(4885);
VN_in_sig(3987)	<=	CN_out_sig(4886);
VN_in_sig(5095)	<=	CN_out_sig(4887);
VN_in_sig(11)	<=	CN_out_sig(4888);
VN_in_sig(787)	<=	CN_out_sig(4889);
VN_in_sig(1511)	<=	CN_out_sig(4890);
VN_in_sig(2151)	<=	CN_out_sig(4891);
VN_in_sig(2847)	<=	CN_out_sig(4892);
VN_in_sig(3575)	<=	CN_out_sig(4893);
VN_in_sig(3991)	<=	CN_out_sig(4894);
VN_in_sig(5099)	<=	CN_out_sig(4895);
VN_in_sig(15)	<=	CN_out_sig(4896);
VN_in_sig(791)	<=	CN_out_sig(4897);
VN_in_sig(1299)	<=	CN_out_sig(4898);
VN_in_sig(2155)	<=	CN_out_sig(4899);
VN_in_sig(2851)	<=	CN_out_sig(4900);
VN_in_sig(3579)	<=	CN_out_sig(4901);
VN_in_sig(3995)	<=	CN_out_sig(4902);
VN_in_sig(5103)	<=	CN_out_sig(4903);
VN_in_sig(19)	<=	CN_out_sig(4904);
VN_in_sig(795)	<=	CN_out_sig(4905);
VN_in_sig(1303)	<=	CN_out_sig(4906);
VN_in_sig(2159)	<=	CN_out_sig(4907);
VN_in_sig(2855)	<=	CN_out_sig(4908);
VN_in_sig(3583)	<=	CN_out_sig(4909);
VN_in_sig(3999)	<=	CN_out_sig(4910);
VN_in_sig(5107)	<=	CN_out_sig(4911);
VN_in_sig(23)	<=	CN_out_sig(4912);
VN_in_sig(799)	<=	CN_out_sig(4913);
VN_in_sig(1307)	<=	CN_out_sig(4914);
VN_in_sig(1947)	<=	CN_out_sig(4915);
VN_in_sig(2859)	<=	CN_out_sig(4916);
VN_in_sig(3587)	<=	CN_out_sig(4917);
VN_in_sig(4003)	<=	CN_out_sig(4918);
VN_in_sig(5111)	<=	CN_out_sig(4919);
VN_in_sig(27)	<=	CN_out_sig(4920);
VN_in_sig(803)	<=	CN_out_sig(4921);
VN_in_sig(1311)	<=	CN_out_sig(4922);
VN_in_sig(1951)	<=	CN_out_sig(4923);
VN_in_sig(2863)	<=	CN_out_sig(4924);
VN_in_sig(3591)	<=	CN_out_sig(4925);
VN_in_sig(4007)	<=	CN_out_sig(4926);
VN_in_sig(5115)	<=	CN_out_sig(4927);
VN_in_sig(31)	<=	CN_out_sig(4928);
VN_in_sig(807)	<=	CN_out_sig(4929);
VN_in_sig(1315)	<=	CN_out_sig(4930);
VN_in_sig(1955)	<=	CN_out_sig(4931);
VN_in_sig(2867)	<=	CN_out_sig(4932);
VN_in_sig(3595)	<=	CN_out_sig(4933);
VN_in_sig(4011)	<=	CN_out_sig(4934);
VN_in_sig(5119)	<=	CN_out_sig(4935);
VN_in_sig(35)	<=	CN_out_sig(4936);
VN_in_sig(811)	<=	CN_out_sig(4937);
VN_in_sig(1319)	<=	CN_out_sig(4938);
VN_in_sig(1959)	<=	CN_out_sig(4939);
VN_in_sig(2871)	<=	CN_out_sig(4940);
VN_in_sig(3599)	<=	CN_out_sig(4941);
VN_in_sig(4015)	<=	CN_out_sig(4942);
VN_in_sig(5123)	<=	CN_out_sig(4943);
VN_in_sig(39)	<=	CN_out_sig(4944);
VN_in_sig(815)	<=	CN_out_sig(4945);
VN_in_sig(1323)	<=	CN_out_sig(4946);
VN_in_sig(1963)	<=	CN_out_sig(4947);
VN_in_sig(2875)	<=	CN_out_sig(4948);
VN_in_sig(3603)	<=	CN_out_sig(4949);
VN_in_sig(4019)	<=	CN_out_sig(4950);
VN_in_sig(5127)	<=	CN_out_sig(4951);
VN_in_sig(43)	<=	CN_out_sig(4952);
VN_in_sig(819)	<=	CN_out_sig(4953);
VN_in_sig(1327)	<=	CN_out_sig(4954);
VN_in_sig(1967)	<=	CN_out_sig(4955);
VN_in_sig(2879)	<=	CN_out_sig(4956);
VN_in_sig(3607)	<=	CN_out_sig(4957);
VN_in_sig(4023)	<=	CN_out_sig(4958);
VN_in_sig(5131)	<=	CN_out_sig(4959);
VN_in_sig(47)	<=	CN_out_sig(4960);
VN_in_sig(823)	<=	CN_out_sig(4961);
VN_in_sig(1331)	<=	CN_out_sig(4962);
VN_in_sig(1971)	<=	CN_out_sig(4963);
VN_in_sig(2883)	<=	CN_out_sig(4964);
VN_in_sig(3611)	<=	CN_out_sig(4965);
VN_in_sig(4027)	<=	CN_out_sig(4966);
VN_in_sig(5135)	<=	CN_out_sig(4967);
VN_in_sig(51)	<=	CN_out_sig(4968);
VN_in_sig(827)	<=	CN_out_sig(4969);
VN_in_sig(1335)	<=	CN_out_sig(4970);
VN_in_sig(1975)	<=	CN_out_sig(4971);
VN_in_sig(2887)	<=	CN_out_sig(4972);
VN_in_sig(3615)	<=	CN_out_sig(4973);
VN_in_sig(4031)	<=	CN_out_sig(4974);
VN_in_sig(5139)	<=	CN_out_sig(4975);
VN_in_sig(55)	<=	CN_out_sig(4976);
VN_in_sig(831)	<=	CN_out_sig(4977);
VN_in_sig(1339)	<=	CN_out_sig(4978);
VN_in_sig(1979)	<=	CN_out_sig(4979);
VN_in_sig(2891)	<=	CN_out_sig(4980);
VN_in_sig(3619)	<=	CN_out_sig(4981);
VN_in_sig(4035)	<=	CN_out_sig(4982);
VN_in_sig(5143)	<=	CN_out_sig(4983);
VN_in_sig(59)	<=	CN_out_sig(4984);
VN_in_sig(835)	<=	CN_out_sig(4985);
VN_in_sig(1343)	<=	CN_out_sig(4986);
VN_in_sig(1983)	<=	CN_out_sig(4987);
VN_in_sig(2895)	<=	CN_out_sig(4988);
VN_in_sig(3623)	<=	CN_out_sig(4989);
VN_in_sig(4039)	<=	CN_out_sig(4990);
VN_in_sig(5147)	<=	CN_out_sig(4991);
VN_in_sig(63)	<=	CN_out_sig(4992);
VN_in_sig(839)	<=	CN_out_sig(4993);
VN_in_sig(1347)	<=	CN_out_sig(4994);
VN_in_sig(1987)	<=	CN_out_sig(4995);
VN_in_sig(2899)	<=	CN_out_sig(4996);
VN_in_sig(3627)	<=	CN_out_sig(4997);
VN_in_sig(4043)	<=	CN_out_sig(4998);
VN_in_sig(5151)	<=	CN_out_sig(4999);
VN_in_sig(67)	<=	CN_out_sig(5000);
VN_in_sig(843)	<=	CN_out_sig(5001);
VN_in_sig(1351)	<=	CN_out_sig(5002);
VN_in_sig(1991)	<=	CN_out_sig(5003);
VN_in_sig(2903)	<=	CN_out_sig(5004);
VN_in_sig(3631)	<=	CN_out_sig(5005);
VN_in_sig(4047)	<=	CN_out_sig(5006);
VN_in_sig(5155)	<=	CN_out_sig(5007);
VN_in_sig(71)	<=	CN_out_sig(5008);
VN_in_sig(847)	<=	CN_out_sig(5009);
VN_in_sig(1355)	<=	CN_out_sig(5010);
VN_in_sig(1995)	<=	CN_out_sig(5011);
VN_in_sig(2907)	<=	CN_out_sig(5012);
VN_in_sig(3635)	<=	CN_out_sig(5013);
VN_in_sig(4051)	<=	CN_out_sig(5014);
VN_in_sig(5159)	<=	CN_out_sig(5015);
VN_in_sig(75)	<=	CN_out_sig(5016);
VN_in_sig(851)	<=	CN_out_sig(5017);
VN_in_sig(1359)	<=	CN_out_sig(5018);
VN_in_sig(1999)	<=	CN_out_sig(5019);
VN_in_sig(2911)	<=	CN_out_sig(5020);
VN_in_sig(3639)	<=	CN_out_sig(5021);
VN_in_sig(4055)	<=	CN_out_sig(5022);
VN_in_sig(5163)	<=	CN_out_sig(5023);
VN_in_sig(79)	<=	CN_out_sig(5024);
VN_in_sig(855)	<=	CN_out_sig(5025);
VN_in_sig(1363)	<=	CN_out_sig(5026);
VN_in_sig(2003)	<=	CN_out_sig(5027);
VN_in_sig(2915)	<=	CN_out_sig(5028);
VN_in_sig(3643)	<=	CN_out_sig(5029);
VN_in_sig(4059)	<=	CN_out_sig(5030);
VN_in_sig(5167)	<=	CN_out_sig(5031);
VN_in_sig(83)	<=	CN_out_sig(5032);
VN_in_sig(859)	<=	CN_out_sig(5033);
VN_in_sig(1367)	<=	CN_out_sig(5034);
VN_in_sig(2007)	<=	CN_out_sig(5035);
VN_in_sig(2919)	<=	CN_out_sig(5036);
VN_in_sig(3647)	<=	CN_out_sig(5037);
VN_in_sig(4063)	<=	CN_out_sig(5038);
VN_in_sig(5171)	<=	CN_out_sig(5039);
VN_in_sig(87)	<=	CN_out_sig(5040);
VN_in_sig(863)	<=	CN_out_sig(5041);
VN_in_sig(1371)	<=	CN_out_sig(5042);
VN_in_sig(2011)	<=	CN_out_sig(5043);
VN_in_sig(2923)	<=	CN_out_sig(5044);
VN_in_sig(3651)	<=	CN_out_sig(5045);
VN_in_sig(4067)	<=	CN_out_sig(5046);
VN_in_sig(5175)	<=	CN_out_sig(5047);
VN_in_sig(91)	<=	CN_out_sig(5048);
VN_in_sig(651)	<=	CN_out_sig(5049);
VN_in_sig(1375)	<=	CN_out_sig(5050);
VN_in_sig(2015)	<=	CN_out_sig(5051);
VN_in_sig(2927)	<=	CN_out_sig(5052);
VN_in_sig(3655)	<=	CN_out_sig(5053);
VN_in_sig(4071)	<=	CN_out_sig(5054);
VN_in_sig(5179)	<=	CN_out_sig(5055);
VN_in_sig(95)	<=	CN_out_sig(5056);
VN_in_sig(655)	<=	CN_out_sig(5057);
VN_in_sig(1379)	<=	CN_out_sig(5058);
VN_in_sig(2019)	<=	CN_out_sig(5059);
VN_in_sig(2931)	<=	CN_out_sig(5060);
VN_in_sig(3659)	<=	CN_out_sig(5061);
VN_in_sig(4075)	<=	CN_out_sig(5062);
VN_in_sig(5183)	<=	CN_out_sig(5063);
VN_in_sig(99)	<=	CN_out_sig(5064);
VN_in_sig(659)	<=	CN_out_sig(5065);
VN_in_sig(1383)	<=	CN_out_sig(5066);
VN_in_sig(2023)	<=	CN_out_sig(5067);
VN_in_sig(2935)	<=	CN_out_sig(5068);
VN_in_sig(3663)	<=	CN_out_sig(5069);
VN_in_sig(4079)	<=	CN_out_sig(5070);
VN_in_sig(4971)	<=	CN_out_sig(5071);
VN_in_sig(103)	<=	CN_out_sig(5072);
VN_in_sig(663)	<=	CN_out_sig(5073);
VN_in_sig(1387)	<=	CN_out_sig(5074);
VN_in_sig(2027)	<=	CN_out_sig(5075);
VN_in_sig(2939)	<=	CN_out_sig(5076);
VN_in_sig(3667)	<=	CN_out_sig(5077);
VN_in_sig(4083)	<=	CN_out_sig(5078);
VN_in_sig(4975)	<=	CN_out_sig(5079);
VN_in_sig(107)	<=	CN_out_sig(5080);
VN_in_sig(667)	<=	CN_out_sig(5081);
VN_in_sig(1391)	<=	CN_out_sig(5082);
VN_in_sig(2031)	<=	CN_out_sig(5083);
VN_in_sig(2943)	<=	CN_out_sig(5084);
VN_in_sig(3671)	<=	CN_out_sig(5085);
VN_in_sig(4087)	<=	CN_out_sig(5086);
VN_in_sig(4979)	<=	CN_out_sig(5087);
VN_in_sig(111)	<=	CN_out_sig(5088);
VN_in_sig(671)	<=	CN_out_sig(5089);
VN_in_sig(1395)	<=	CN_out_sig(5090);
VN_in_sig(2035)	<=	CN_out_sig(5091);
VN_in_sig(2947)	<=	CN_out_sig(5092);
VN_in_sig(3459)	<=	CN_out_sig(5093);
VN_in_sig(4091)	<=	CN_out_sig(5094);
VN_in_sig(4983)	<=	CN_out_sig(5095);
VN_in_sig(115)	<=	CN_out_sig(5096);
VN_in_sig(675)	<=	CN_out_sig(5097);
VN_in_sig(1399)	<=	CN_out_sig(5098);
VN_in_sig(2039)	<=	CN_out_sig(5099);
VN_in_sig(2951)	<=	CN_out_sig(5100);
VN_in_sig(3463)	<=	CN_out_sig(5101);
VN_in_sig(4095)	<=	CN_out_sig(5102);
VN_in_sig(4987)	<=	CN_out_sig(5103);
VN_in_sig(119)	<=	CN_out_sig(5104);
VN_in_sig(679)	<=	CN_out_sig(5105);
VN_in_sig(1403)	<=	CN_out_sig(5106);
VN_in_sig(2043)	<=	CN_out_sig(5107);
VN_in_sig(2955)	<=	CN_out_sig(5108);
VN_in_sig(3467)	<=	CN_out_sig(5109);
VN_in_sig(4099)	<=	CN_out_sig(5110);
VN_in_sig(4991)	<=	CN_out_sig(5111);
VN_in_sig(123)	<=	CN_out_sig(5112);
VN_in_sig(683)	<=	CN_out_sig(5113);
VN_in_sig(1407)	<=	CN_out_sig(5114);
VN_in_sig(2047)	<=	CN_out_sig(5115);
VN_in_sig(2959)	<=	CN_out_sig(5116);
VN_in_sig(3471)	<=	CN_out_sig(5117);
VN_in_sig(4103)	<=	CN_out_sig(5118);
VN_in_sig(4995)	<=	CN_out_sig(5119);
VN_in_sig(127)	<=	CN_out_sig(5120);
VN_in_sig(687)	<=	CN_out_sig(5121);
VN_in_sig(1411)	<=	CN_out_sig(5122);
VN_in_sig(2051)	<=	CN_out_sig(5123);
VN_in_sig(2963)	<=	CN_out_sig(5124);
VN_in_sig(3475)	<=	CN_out_sig(5125);
VN_in_sig(3891)	<=	CN_out_sig(5126);
VN_in_sig(4999)	<=	CN_out_sig(5127);
VN_in_sig(131)	<=	CN_out_sig(5128);
VN_in_sig(691)	<=	CN_out_sig(5129);
VN_in_sig(1415)	<=	CN_out_sig(5130);
VN_in_sig(2055)	<=	CN_out_sig(5131);
VN_in_sig(2967)	<=	CN_out_sig(5132);
VN_in_sig(3479)	<=	CN_out_sig(5133);
VN_in_sig(3895)	<=	CN_out_sig(5134);
VN_in_sig(5003)	<=	CN_out_sig(5135);
VN_in_sig(135)	<=	CN_out_sig(5136);
VN_in_sig(695)	<=	CN_out_sig(5137);
VN_in_sig(1419)	<=	CN_out_sig(5138);
VN_in_sig(2059)	<=	CN_out_sig(5139);
VN_in_sig(2971)	<=	CN_out_sig(5140);
VN_in_sig(3483)	<=	CN_out_sig(5141);
VN_in_sig(3899)	<=	CN_out_sig(5142);
VN_in_sig(5007)	<=	CN_out_sig(5143);
VN_in_sig(139)	<=	CN_out_sig(5144);
VN_in_sig(699)	<=	CN_out_sig(5145);
VN_in_sig(1423)	<=	CN_out_sig(5146);
VN_in_sig(2063)	<=	CN_out_sig(5147);
VN_in_sig(2975)	<=	CN_out_sig(5148);
VN_in_sig(3487)	<=	CN_out_sig(5149);
VN_in_sig(3903)	<=	CN_out_sig(5150);
VN_in_sig(5011)	<=	CN_out_sig(5151);
VN_in_sig(143)	<=	CN_out_sig(5152);
VN_in_sig(703)	<=	CN_out_sig(5153);
VN_in_sig(1427)	<=	CN_out_sig(5154);
VN_in_sig(2067)	<=	CN_out_sig(5155);
VN_in_sig(2979)	<=	CN_out_sig(5156);
VN_in_sig(3491)	<=	CN_out_sig(5157);
VN_in_sig(3907)	<=	CN_out_sig(5158);
VN_in_sig(5015)	<=	CN_out_sig(5159);
VN_in_sig(147)	<=	CN_out_sig(5160);
VN_in_sig(707)	<=	CN_out_sig(5161);
VN_in_sig(1431)	<=	CN_out_sig(5162);
VN_in_sig(2071)	<=	CN_out_sig(5163);
VN_in_sig(2983)	<=	CN_out_sig(5164);
VN_in_sig(3495)	<=	CN_out_sig(5165);
VN_in_sig(3911)	<=	CN_out_sig(5166);
VN_in_sig(5019)	<=	CN_out_sig(5167);
VN_in_sig(151)	<=	CN_out_sig(5168);
VN_in_sig(711)	<=	CN_out_sig(5169);
VN_in_sig(1435)	<=	CN_out_sig(5170);
VN_in_sig(2075)	<=	CN_out_sig(5171);
VN_in_sig(2987)	<=	CN_out_sig(5172);
VN_in_sig(3499)	<=	CN_out_sig(5173);
VN_in_sig(3915)	<=	CN_out_sig(5174);
VN_in_sig(5023)	<=	CN_out_sig(5175);
VN_in_sig(155)	<=	CN_out_sig(5176);
VN_in_sig(715)	<=	CN_out_sig(5177);
VN_in_sig(1439)	<=	CN_out_sig(5178);
VN_in_sig(2079)	<=	CN_out_sig(5179);
VN_in_sig(2991)	<=	CN_out_sig(5180);
VN_in_sig(3503)	<=	CN_out_sig(5181);
VN_in_sig(3919)	<=	CN_out_sig(5182);
VN_in_sig(5027)	<=	CN_out_sig(5183);


