----------------------------------------------------------------------------------
-- Engineer: Burak UNAL 
-- 
-- Create Date:    
-- Design Name:  Created by Burak UNAL 
-- Project Name: Gallager-B Hard decision Bit-Flipping algorithm
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--COPYRIGHT            : burak@email.arizona.edu
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE ieee.std_logic_unsigned.all;

entity random_numb is
    generic ( width : integer :=  31;
              threshold : integer:= 1717986918	 );
port (
      clk, ena : in std_logic;
		
      ran_out  		: out STD_LOGIC_VECTOR(1295 downto 0)
    );
end random_numb;

architecture Behavioral of random_numb is
signal tempo        : std_logic_vector(width-1 downto 0);
signal ran_out_sig  : STD_LOGIC_VECTOR(1295 downto 0):="000001100001000000000010000010000100000000100000100000100000100001000010000000010010010001000010000010000010000100000010000100000100000000001100000010000000100000100000000100000001000000000100000001000000000010000100001000000100000011000010100100101110010010100010001001000010010010000100100100101010100011010100010001001010101010001001001010001010101000010010010000100100010001100101000001000101000001001001000001010010000010100100000110000100001111000011000010000001000100001000010010001000000101000001000001000100000100001000001000000000010000001000000100000000100000010000100100000001000000000001000000000001000000000001000000000000100000000000001000000000000000100000000000000000010000000000000010000000000000000100000000000000100000000000000000100000000000000001000000000000000000100000000000000001000000000000000001000000000000100000000000000010000000000000100000000000000010000000000001000000000000100111000000100111100011100001001000010000100000001100000000100001111000001000000011100001000000011100000010100000011100010000001110000100000011100000100001110000011100100000110001100001000001001000111000000100100001010000100100000010001001100010011100000100010000100001000010011100001000010010010010000010000000100010000010000010010001000000100010000100010000000100100010000100001000000011";

begin
process(clk)
variable rand_temp : std_logic_vector(width-1 downto 0):="110"& X"1254EA7"; 
variable temp : std_logic := '0';
begin
	if(rising_edge(clk) and ena='1') then
	temp := rand_temp(width-1) xor rand_temp(width-2);
	rand_temp(width-1 downto 1) := rand_temp(width-2 downto 0);
	rand_temp(0) := temp;
	
	ran_out_sig(1295 downto 1) <= ran_out_sig(1294 downto 0);
			if (rand_temp < threshold) then
			ran_out_sig(0) <= '0';
	       else
			ran_out_sig (0) <='1';
			end if;
			
	 
	end if;

	
end process;
ran_out <= ran_out_sig;
end;
