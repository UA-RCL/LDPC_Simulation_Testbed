 ----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity encoder is
    Port ( 	clk			: in	STD_LOGIC;
			rst			: in	STD_LOGIC;
			init		: in	STD_LOGIC;
			start		: in	STD_LOGIC;
			threshold	:in std_logic_vector(14 downto 0);

		
            codeword_out	: out std_logic_vector(99 downto 0);
			codeword_avail	: out	STD_LOGIC);
end encoder;

architecture rtl of encoder is
COMPONENT reg_unit is
    Port ( clk			: in	STD_LOGIC;
			rst			: in	STD_LOGIC;
			init		: in	STD_LOGIC;
			start		: in	STD_LOGIC;
			data_init	: in std_logic_vector(149 downto 0);
			threshold	: in std_logic_vector(14 downto 0);         
           
           ran_bit			: out	STD_LOGIC);
end COMPONENT;

signal codeword_out_sig: 	std_logic_vector (99 downto 0);

signal   reg_sig_0:     std_logic_vector (149 downto 0);
signal   reg_sig_1:     std_logic_vector (149 downto 0);
signal   reg_sig_2:     std_logic_vector (149 downto 0);
signal   reg_sig_3:     std_logic_vector (149 downto 0);
signal   reg_sig_4:     std_logic_vector (149 downto 0);
signal   reg_sig_5:     std_logic_vector (149 downto 0);
signal   reg_sig_6:     std_logic_vector (149 downto 0);
signal   reg_sig_7:     std_logic_vector (149 downto 0);
signal   reg_sig_8:     std_logic_vector (149 downto 0);
signal   reg_sig_9:     std_logic_vector (149 downto 0);
signal   reg_sig_10:    std_logic_vector (149 downto 0);
signal   reg_sig_11:    std_logic_vector (149 downto 0);
signal   reg_sig_12:    std_logic_vector (149 downto 0);
signal   reg_sig_13:    std_logic_vector (149 downto 0);
signal   reg_sig_14:    std_logic_vector (149 downto 0);
signal   reg_sig_15:    std_logic_vector (149 downto 0);
signal   reg_sig_16:    std_logic_vector (149 downto 0);
signal   reg_sig_17:    std_logic_vector (149 downto 0);
signal   reg_sig_18:    std_logic_vector (149 downto 0);
signal   reg_sig_19:    std_logic_vector (149 downto 0);
signal   reg_sig_20:    std_logic_vector (149 downto 0);
signal   reg_sig_21:    std_logic_vector (149 downto 0);
signal   reg_sig_22:    std_logic_vector (149 downto 0);
signal   reg_sig_23:    std_logic_vector (149 downto 0);
signal   reg_sig_24:    std_logic_vector (149 downto 0);
signal   reg_sig_25:    std_logic_vector (149 downto 0);
signal   reg_sig_26:    std_logic_vector (149 downto 0);
signal   reg_sig_27:    std_logic_vector (149 downto 0);
signal   reg_sig_28:    std_logic_vector (149 downto 0);
signal   reg_sig_29:    std_logic_vector (149 downto 0);
signal   reg_sig_30:    std_logic_vector (149 downto 0);
signal   reg_sig_31:    std_logic_vector (149 downto 0);
signal   reg_sig_32:    std_logic_vector (149 downto 0);
signal   reg_sig_33:    std_logic_vector (149 downto 0);
signal   reg_sig_34:    std_logic_vector (149 downto 0);
signal   reg_sig_35:    std_logic_vector (149 downto 0);
signal   reg_sig_36:    std_logic_vector (149 downto 0);
signal   reg_sig_37:    std_logic_vector (149 downto 0);
signal   reg_sig_38:    std_logic_vector (149 downto 0);
signal   reg_sig_39:    std_logic_vector (149 downto 0);
signal   reg_sig_40:    std_logic_vector (149 downto 0);
signal   reg_sig_41:    std_logic_vector (149 downto 0);
signal   reg_sig_42:    std_logic_vector (149 downto 0);
signal   reg_sig_43:    std_logic_vector (149 downto 0);
signal   reg_sig_44:    std_logic_vector (149 downto 0);
signal   reg_sig_45:    std_logic_vector (149 downto 0);
signal   reg_sig_46:    std_logic_vector (149 downto 0);
signal   reg_sig_47:    std_logic_vector (149 downto 0);
signal   reg_sig_48:    std_logic_vector (149 downto 0);
signal   reg_sig_49:    std_logic_vector (149 downto 0);
signal   reg_sig_50:    std_logic_vector (149 downto 0);
signal   reg_sig_51:    std_logic_vector (149 downto 0);
signal   reg_sig_52:    std_logic_vector (149 downto 0);
signal   reg_sig_53:    std_logic_vector (149 downto 0);
signal   reg_sig_54:    std_logic_vector (149 downto 0);
signal   reg_sig_55:    std_logic_vector (149 downto 0);
signal   reg_sig_56:    std_logic_vector (149 downto 0);
signal   reg_sig_57:    std_logic_vector (149 downto 0);
signal   reg_sig_58:    std_logic_vector (149 downto 0);
signal   reg_sig_59:    std_logic_vector (149 downto 0);
signal   reg_sig_60:    std_logic_vector (149 downto 0);
signal   reg_sig_61:    std_logic_vector (149 downto 0);
signal   reg_sig_62:    std_logic_vector (149 downto 0);
signal   reg_sig_63:    std_logic_vector (149 downto 0);
signal   reg_sig_64:    std_logic_vector (149 downto 0);
signal   reg_sig_65:    std_logic_vector (149 downto 0);
signal   reg_sig_66:    std_logic_vector (149 downto 0);
signal   reg_sig_67:    std_logic_vector (149 downto 0);
signal   reg_sig_68:    std_logic_vector (149 downto 0);
signal   reg_sig_69:    std_logic_vector (149 downto 0);
signal   reg_sig_70:    std_logic_vector (149 downto 0);
signal   reg_sig_71:    std_logic_vector (149 downto 0);
signal   reg_sig_72:    std_logic_vector (149 downto 0);
signal   reg_sig_73:    std_logic_vector (149 downto 0);
signal   reg_sig_74:    std_logic_vector (149 downto 0);
signal   reg_sig_75:    std_logic_vector (149 downto 0);
signal   reg_sig_76:    std_logic_vector (149 downto 0);
signal   reg_sig_77:    std_logic_vector (149 downto 0);
signal   reg_sig_78:    std_logic_vector (149 downto 0);
signal   reg_sig_79:    std_logic_vector (149 downto 0);
signal   reg_sig_80:    std_logic_vector (149 downto 0);
signal   reg_sig_81:    std_logic_vector (149 downto 0);
signal   reg_sig_82:    std_logic_vector (149 downto 0);
signal   reg_sig_83:    std_logic_vector (149 downto 0);
signal   reg_sig_84:    std_logic_vector (149 downto 0);
signal   reg_sig_85:    std_logic_vector (149 downto 0);
signal   reg_sig_86:    std_logic_vector (149 downto 0);
signal   reg_sig_87:    std_logic_vector (149 downto 0);
signal   reg_sig_88:    std_logic_vector (149 downto 0);
signal   reg_sig_89:    std_logic_vector (149 downto 0);
signal   reg_sig_90:    std_logic_vector (149 downto 0);
signal   reg_sig_91:    std_logic_vector (149 downto 0);
signal   reg_sig_92:    std_logic_vector (149 downto 0);
signal   reg_sig_93:    std_logic_vector (149 downto 0);
signal   reg_sig_94:    std_logic_vector (149 downto 0);
signal   reg_sig_95:    std_logic_vector (149 downto 0);
signal   reg_sig_96:    std_logic_vector (149 downto 0);
signal   reg_sig_97:    std_logic_vector (149 downto 0);
signal   reg_sig_98:    std_logic_vector (149 downto 0);
signal   reg_sig_99:    std_logic_vector (149 downto 0);


begin

reg_unit_0     : reg_unit port map (clk, rst, init, start, reg_sig_0,threshold,codeword_out_sig(0));
reg_unit_1     : reg_unit port map (clk, rst, init, start, reg_sig_1,threshold,codeword_out_sig(1));
reg_unit_2     : reg_unit port map (clk, rst, init, start, reg_sig_2,threshold,codeword_out_sig(2));
reg_unit_3     : reg_unit port map (clk, rst, init, start, reg_sig_3,threshold,codeword_out_sig(3));
reg_unit_4     : reg_unit port map (clk, rst, init, start, reg_sig_4,threshold,codeword_out_sig(4));
reg_unit_5     : reg_unit port map (clk, rst, init, start, reg_sig_5,threshold,codeword_out_sig(5));
reg_unit_6     : reg_unit port map (clk, rst, init, start, reg_sig_6,threshold,codeword_out_sig(6));
reg_unit_7     : reg_unit port map (clk, rst, init, start, reg_sig_7,threshold,codeword_out_sig(7));
reg_unit_8     : reg_unit port map (clk, rst, init, start, reg_sig_8,threshold,codeword_out_sig(8));
reg_unit_9     : reg_unit port map (clk, rst, init, start, reg_sig_9,threshold,codeword_out_sig(9));
reg_unit_10    : reg_unit port map (clk, rst, init, start, reg_sig_10,threshold,codeword_out_sig(10));
reg_unit_11    : reg_unit port map (clk, rst, init, start, reg_sig_11,threshold,codeword_out_sig(11));
reg_unit_12    : reg_unit port map (clk, rst, init, start, reg_sig_12,threshold,codeword_out_sig(12));
reg_unit_13    : reg_unit port map (clk, rst, init, start, reg_sig_13,threshold,codeword_out_sig(13));
reg_unit_14    : reg_unit port map (clk, rst, init, start, reg_sig_14,threshold,codeword_out_sig(14));
reg_unit_15    : reg_unit port map (clk, rst, init, start, reg_sig_15,threshold,codeword_out_sig(15));
reg_unit_16    : reg_unit port map (clk, rst, init, start, reg_sig_16,threshold,codeword_out_sig(16));
reg_unit_17    : reg_unit port map (clk, rst, init, start, reg_sig_17,threshold,codeword_out_sig(17));
reg_unit_18    : reg_unit port map (clk, rst, init, start, reg_sig_18,threshold,codeword_out_sig(18));
reg_unit_19    : reg_unit port map (clk, rst, init, start, reg_sig_19,threshold,codeword_out_sig(19));
reg_unit_20    : reg_unit port map (clk, rst, init, start, reg_sig_20,threshold,codeword_out_sig(20));
reg_unit_21    : reg_unit port map (clk, rst, init, start, reg_sig_21,threshold,codeword_out_sig(21));
reg_unit_22    : reg_unit port map (clk, rst, init, start, reg_sig_22,threshold,codeword_out_sig(22));
reg_unit_23    : reg_unit port map (clk, rst, init, start, reg_sig_23,threshold,codeword_out_sig(23));
reg_unit_24    : reg_unit port map (clk, rst, init, start, reg_sig_24,threshold,codeword_out_sig(24));
reg_unit_25    : reg_unit port map (clk, rst, init, start, reg_sig_25,threshold,codeword_out_sig(25));
reg_unit_26    : reg_unit port map (clk, rst, init, start, reg_sig_26,threshold,codeword_out_sig(26));
reg_unit_27    : reg_unit port map (clk, rst, init, start, reg_sig_27,threshold,codeword_out_sig(27));
reg_unit_28    : reg_unit port map (clk, rst, init, start, reg_sig_28,threshold,codeword_out_sig(28));
reg_unit_29    : reg_unit port map (clk, rst, init, start, reg_sig_29,threshold,codeword_out_sig(29));
reg_unit_30    : reg_unit port map (clk, rst, init, start, reg_sig_30,threshold,codeword_out_sig(30));
reg_unit_31    : reg_unit port map (clk, rst, init, start, reg_sig_31,threshold,codeword_out_sig(31));
reg_unit_32    : reg_unit port map (clk, rst, init, start, reg_sig_32,threshold,codeword_out_sig(32));
reg_unit_33    : reg_unit port map (clk, rst, init, start, reg_sig_33,threshold,codeword_out_sig(33));
reg_unit_34    : reg_unit port map (clk, rst, init, start, reg_sig_34,threshold,codeword_out_sig(34));
reg_unit_35    : reg_unit port map (clk, rst, init, start, reg_sig_35,threshold,codeword_out_sig(35));
reg_unit_36    : reg_unit port map (clk, rst, init, start, reg_sig_36,threshold,codeword_out_sig(36));
reg_unit_37    : reg_unit port map (clk, rst, init, start, reg_sig_37,threshold,codeword_out_sig(37));
reg_unit_38    : reg_unit port map (clk, rst, init, start, reg_sig_38,threshold,codeword_out_sig(38));
reg_unit_39    : reg_unit port map (clk, rst, init, start, reg_sig_39,threshold,codeword_out_sig(39));
reg_unit_40    : reg_unit port map (clk, rst, init, start, reg_sig_40,threshold,codeword_out_sig(40));
reg_unit_41    : reg_unit port map (clk, rst, init, start, reg_sig_41,threshold,codeword_out_sig(41));
reg_unit_42    : reg_unit port map (clk, rst, init, start, reg_sig_42,threshold,codeword_out_sig(42));
reg_unit_43    : reg_unit port map (clk, rst, init, start, reg_sig_43,threshold,codeword_out_sig(43));
reg_unit_44    : reg_unit port map (clk, rst, init, start, reg_sig_44,threshold,codeword_out_sig(44));
reg_unit_45    : reg_unit port map (clk, rst, init, start, reg_sig_45,threshold,codeword_out_sig(45));
reg_unit_46    : reg_unit port map (clk, rst, init, start, reg_sig_46,threshold,codeword_out_sig(46));
reg_unit_47    : reg_unit port map (clk, rst, init, start, reg_sig_47,threshold,codeword_out_sig(47));
reg_unit_48    : reg_unit port map (clk, rst, init, start, reg_sig_48,threshold,codeword_out_sig(48));
reg_unit_49    : reg_unit port map (clk, rst, init, start, reg_sig_49,threshold,codeword_out_sig(49));
reg_unit_50    : reg_unit port map (clk, rst, init, start, reg_sig_50,threshold,codeword_out_sig(50));
reg_unit_51    : reg_unit port map (clk, rst, init, start, reg_sig_51,threshold,codeword_out_sig(51));
reg_unit_52    : reg_unit port map (clk, rst, init, start, reg_sig_52,threshold,codeword_out_sig(52));
reg_unit_53    : reg_unit port map (clk, rst, init, start, reg_sig_53,threshold,codeword_out_sig(53));
reg_unit_54    : reg_unit port map (clk, rst, init, start, reg_sig_54,threshold,codeword_out_sig(54));
reg_unit_55    : reg_unit port map (clk, rst, init, start, reg_sig_55,threshold,codeword_out_sig(55));
reg_unit_56    : reg_unit port map (clk, rst, init, start, reg_sig_56,threshold,codeword_out_sig(56));
reg_unit_57    : reg_unit port map (clk, rst, init, start, reg_sig_57,threshold,codeword_out_sig(57));
reg_unit_58    : reg_unit port map (clk, rst, init, start, reg_sig_58,threshold,codeword_out_sig(58));
reg_unit_59    : reg_unit port map (clk, rst, init, start, reg_sig_59,threshold,codeword_out_sig(59));
reg_unit_60    : reg_unit port map (clk, rst, init, start, reg_sig_60,threshold,codeword_out_sig(60));
reg_unit_61    : reg_unit port map (clk, rst, init, start, reg_sig_61,threshold,codeword_out_sig(61));
reg_unit_62    : reg_unit port map (clk, rst, init, start, reg_sig_62,threshold,codeword_out_sig(62));
reg_unit_63    : reg_unit port map (clk, rst, init, start, reg_sig_63,threshold,codeword_out_sig(63));
reg_unit_64    : reg_unit port map (clk, rst, init, start, reg_sig_64,threshold,codeword_out_sig(64));
reg_unit_65    : reg_unit port map (clk, rst, init, start, reg_sig_65,threshold,codeword_out_sig(65));
reg_unit_66    : reg_unit port map (clk, rst, init, start, reg_sig_66,threshold,codeword_out_sig(66));
reg_unit_67    : reg_unit port map (clk, rst, init, start, reg_sig_67,threshold,codeword_out_sig(67));
reg_unit_68    : reg_unit port map (clk, rst, init, start, reg_sig_68,threshold,codeword_out_sig(68));
reg_unit_69    : reg_unit port map (clk, rst, init, start, reg_sig_69,threshold,codeword_out_sig(69));
reg_unit_70    : reg_unit port map (clk, rst, init, start, reg_sig_70,threshold,codeword_out_sig(70));
reg_unit_71    : reg_unit port map (clk, rst, init, start, reg_sig_71,threshold,codeword_out_sig(71));
reg_unit_72    : reg_unit port map (clk, rst, init, start, reg_sig_72,threshold,codeword_out_sig(72));
reg_unit_73    : reg_unit port map (clk, rst, init, start, reg_sig_73,threshold,codeword_out_sig(73));
reg_unit_74    : reg_unit port map (clk, rst, init, start, reg_sig_74,threshold,codeword_out_sig(74));
reg_unit_75    : reg_unit port map (clk, rst, init, start, reg_sig_75,threshold,codeword_out_sig(75));
reg_unit_76    : reg_unit port map (clk, rst, init, start, reg_sig_76,threshold,codeword_out_sig(76));
reg_unit_77    : reg_unit port map (clk, rst, init, start, reg_sig_77,threshold,codeword_out_sig(77));
reg_unit_78    : reg_unit port map (clk, rst, init, start, reg_sig_78,threshold,codeword_out_sig(78));
reg_unit_79    : reg_unit port map (clk, rst, init, start, reg_sig_79,threshold,codeword_out_sig(79));
reg_unit_80    : reg_unit port map (clk, rst, init, start, reg_sig_80,threshold,codeword_out_sig(80));
reg_unit_81    : reg_unit port map (clk, rst, init, start, reg_sig_81,threshold,codeword_out_sig(81));
reg_unit_82    : reg_unit port map (clk, rst, init, start, reg_sig_82,threshold,codeword_out_sig(82));
reg_unit_83    : reg_unit port map (clk, rst, init, start, reg_sig_83,threshold,codeword_out_sig(83));
reg_unit_84    : reg_unit port map (clk, rst, init, start, reg_sig_84,threshold,codeword_out_sig(84));
reg_unit_85    : reg_unit port map (clk, rst, init, start, reg_sig_85,threshold,codeword_out_sig(85));
reg_unit_86    : reg_unit port map (clk, rst, init, start, reg_sig_86,threshold,codeword_out_sig(86));
reg_unit_87    : reg_unit port map (clk, rst, init, start, reg_sig_87,threshold,codeword_out_sig(87));
reg_unit_88    : reg_unit port map (clk, rst, init, start, reg_sig_88,threshold,codeword_out_sig(88));
reg_unit_89    : reg_unit port map (clk, rst, init, start, reg_sig_89,threshold,codeword_out_sig(89));
reg_unit_90    : reg_unit port map (clk, rst, init, start, reg_sig_90,threshold,codeword_out_sig(90));
reg_unit_91    : reg_unit port map (clk, rst, init, start, reg_sig_91,threshold,codeword_out_sig(91));
reg_unit_92    : reg_unit port map (clk, rst, init, start, reg_sig_92,threshold,codeword_out_sig(92));
reg_unit_93    : reg_unit port map (clk, rst, init, start, reg_sig_93,threshold,codeword_out_sig(93));
reg_unit_94    : reg_unit port map (clk, rst, init, start, reg_sig_94,threshold,codeword_out_sig(94));
reg_unit_95    : reg_unit port map (clk, rst, init, start, reg_sig_95,threshold,codeword_out_sig(95));
reg_unit_96    : reg_unit port map (clk, rst, init, start, reg_sig_96,threshold,codeword_out_sig(96));
reg_unit_97    : reg_unit port map (clk, rst, init, start, reg_sig_97,threshold,codeword_out_sig(97));
reg_unit_98    : reg_unit port map (clk, rst, init, start, reg_sig_98,threshold,codeword_out_sig(98));
reg_unit_99    : reg_unit port map (clk, rst, init, start, reg_sig_99,threshold,codeword_out_sig(99));

codeword_out <= codeword_out_sig;

process(clk)
begin
	if clk'event and clk = '1' then
		if rst = '1' then
reg_sig_0       <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_1       <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_2       <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_3       <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_4       <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_5       <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_6       <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_7       <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_8       <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_9       <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_10      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_11      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_12      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_13      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_14      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_15      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_16      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_17      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_18      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_19      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_20      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_21      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_22      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_23      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_24      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_25      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_26      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_27      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_28      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_29      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_30      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_31      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_32      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_33      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_34      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_35      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_36      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_37      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_38      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_39      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_40      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_41      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_42      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_43      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_44      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_45      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_46      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_47      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_48      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_49      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_50      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_51      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_52      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_53      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_54      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_55      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_56      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_57      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_58      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_59      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_60      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_61      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_62      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_63      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_64      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_65      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_66      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_67      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_68      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_69      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_70      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_71      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_72      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_73      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_74      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_75      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_76      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_77      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_78      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_79      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_80      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_81      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_82      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_83      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_84      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_85      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_86      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_87      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_88      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_89      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_90      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_91      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_92      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_93      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_94      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_95      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_96      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_97      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_98      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
reg_sig_99      <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

		elsif init='1' then
reg_sig_0       <= "110100101000110000100110110000000010011011111000101100001011010010110111011011001001100001001011011110100000100001101010100100001110011010100110101110";
reg_sig_1       <= "110110011111100011111100101110000000000010111001010011010100000111010111111010010101011000011111001100011010100101011100011110111010001010001000101010";
reg_sig_2       <= "011011110000100111101111011101011101100100100101110111000001110110001000101110000111000100010100001101001110000111001101111111110110110110110100010101";
reg_sig_3       <= "010011001101000100100010011010101111010100111101111111001101001011101110001111010101001010100100010101101010100101001001001100011010111001100100101101";
reg_sig_4       <= "100010011110100000111100010111011001011100011100110001000110101111001111101100001001011010010101101010100001010001100011011110011110010111001100100010";
reg_sig_5       <= "111111111110001010010010100101100001011011010111001000110100110110100110101110110110110011110001001010011100100101100100000011111101010100111011111100";
reg_sig_6       <= "010100010000000000100110111101100001111001000010011110111110011100101000111011001001010101001000101111100111111011010011101110011010000110100100011101";
reg_sig_7       <= "011010101000100001001011010100000101001000000011001011001101001011100010000000001100110011010110101000110011100100110011110010010100010001100111111011";
reg_sig_8       <= "011011100111100010001110011111101001111011101111110000111101111111111110101011000110111000010000011101110001001011111101011111010000011000011110100001";
reg_sig_9       <= "100110111101111011100111001110101110111010011011000011011011111011110011101101000001111101110011101010110101010011111000111000101010111010010011100110";
reg_sig_10      <= "110010111101110100100011101101000100000111110110101111101110011101010111111100011010000101110011011011111001111100001000110110100100010101111100110101";
reg_sig_11      <= "010000010001111001100110110000110101100101010001100101110111100010011100101111011000100110001000011011101101001011001011111110100101101111011100001110";
reg_sig_12      <= "010101110000010000011010101000100110110011111111100000011111111110101111011001000000100000111010110110100101010011001111110100110011010111011111001001";
reg_sig_13      <= "011110010111110100001011101010101111111110001110111110010011010101110000010001110001011101100010100101000010001011110100010000111010001100100101101110";
reg_sig_14      <= "000011101011110010011011001101110011000001010100111100000110011000001011001100111111111110110100101001111001101111010101101110011001111010101101100111";
reg_sig_15      <= "010111100110100110000110101100000111100010001000100000001111010011010010010101110111011001011010011101010100010011110111100111001110000111111001000011";
reg_sig_16      <= "100100111100101111111111100101111001111000011100100000110110111110100111110011000000100000010010000100101110010000000011010110011010111001010000010011";
reg_sig_17      <= "111001110100010111101100001001100110000000001110110110010111010000011110000111000010110100100100000001100011001010011000010011011101011000001100110110";
reg_sig_18      <= "110011001000111010000010011000100001110100010011101110100101000101001100000101010110100101010001010000010000110001101110011011111010101011011001111011";
reg_sig_19      <= "110110001011111100110000001101100011101111000100001011101101110001011110011001000001101011100110000000101100000001100011011001110111111100110101100101";
reg_sig_20      <= "100010000010001010110000110110010011111100111101011011110011100010111110011010100101001110001100010100001011100011111001111110001101011110111011101001";
reg_sig_21      <= "001001101101100110000101001111111001011010011000000011101110110111110100111101011100001000001001010110010001111101010001011110111010011001100101010010";
reg_sig_22      <= "001010011100101001101010111010110111011110101001010010110100001110101100100001110001000111100101111010000011110111100010100000110100000101010110010110";
reg_sig_23      <= "101001100011110011101011010011010101101011001000000110100010100001010111001010001001000000110011000011110011100000001111011101100001000101100011011001";
reg_sig_24      <= "011110100000101110000010101011101111100110110010100010011110001010101110000010000011000010001111010111111101101000001110100100100000011011011110100111";
reg_sig_25      <= "111001010011100001001000011100001101000100100011100001100011101000111001111101110011010100101001111000110010111100010010110001000001110101100111000010";
reg_sig_26      <= "101100100111110110010000010111000110000111001101111011011010100001010001110011010011000110111100010010110001110001010001010111111010001111100101100110";
reg_sig_27      <= "110010001011101100100001101100000111001010111110011111111101100110001011001001111000111011011101011000100011101010101111100101010000011000010001010001";
reg_sig_28      <= "100111100000010001001001110100111000001111001000000101011111001001111110101111010000010000001110000111011001000111110101010110010011000111011111101101";
reg_sig_29      <= "110101011101010111010101110011101011000001001001001011011001011101111111001001011000100011001111001111011100010011111111110010001110101001011111001111";
reg_sig_30      <= "001001111011101101010100011111110110111010101100100000111011001101000111110000010111101011100011011010000010100111010000001001011010100110100111001011";
reg_sig_31      <= "010000111010111000001010001000111000011111111101001000111010111000110011111010010110111100111100010101101111001101101101011000011010110111111100101001";
reg_sig_32      <= "001100111011011101010001000101110111001110111001111000111011001110010101101110100011110101110110011111100100100111100110001101110100101101001110001100";
reg_sig_33      <= "100101100111110110100000101001111001011110001101100000001001111000110101111101110111010111100000010110101010110111100000111111110010101111110001000100";
reg_sig_34      <= "111110100011100100011110011011001010111011011010010110111101010100000100001111001001000111001001111011100011011000110011001100001111000111000100001110";
reg_sig_35      <= "000110100111101111101110010011010101011111011110110000010010100011110001101000110100001101110110001111101111111000101110101110110101011010000100101001";
reg_sig_36      <= "000101001010100001111100100111010101010111010011110011111110100001110110101111010011100100000010100110001100100101010010100000100011101001110000111001";
reg_sig_37      <= "100100100010111010000110111010101101100001000001010001011011011011110100111000001101000111011010011000111101110101000110001010110000101001001000011100";
reg_sig_38      <= "110000101101011001110111111100110101000100010101011011101010011011100100100110011000000101111011101011011101010110100010100001001000100010011010010101";
reg_sig_39      <= "100010011101111011010100001010111001110001101111001000000001001110011011110001111001110111111111000011000011011000011110001100100010111100000011111100";
reg_sig_40      <= "100110101111000001101111000100100011001011000010110010111000010001100110000010111101000010111100000101010101000111101101110001011001100100100010001011";
reg_sig_41      <= "100010000100110111101111101110100111011000101110000010000101101100010011101000000110001000101001111011011000010101000101110110001011110100111110011011";
reg_sig_42      <= "000100010001111011001101101110110101110110111101000100111101111010011101011001010100101011011100100111010111100011001100101000101100110010001111011111";
reg_sig_43      <= "100100111100100110011000100111110001100000111100111001001011101000100001101111001001010100100101001011100001001101111010110100110110011010111011000100";
reg_sig_44      <= "111010011111010010100010100010001100110100011000110001000100111011001110000111101101001100011010000011001001101000101011100011001000111010111111111011";
reg_sig_45      <= "100001100001000110010000010011100010011010010111010111100111111100011011100110101001000110010100000101101011001011010110000100111011111101110111010001";
reg_sig_46      <= "011100011011000111101110011001001011101111011001010001001001000011010101101101011010011010011010011100001000011001110101001100100001101011111000010111";
reg_sig_47      <= "110010101110110100100011101111101111101001001010110100011010011011100111110101001111100010110100101001000111011001100000010001010100111101001101011010";
reg_sig_48      <= "011111001110110110000110111001000100110111011001111010111100111000000111010101010111000011110111011011001101011011110111000110001010011000100000110111";
reg_sig_49      <= "101001001000000100110000101001001101011101010101010100101110010010010001001000000000110000110111110100000011101010001000100001001101011110101010011011";
reg_sig_50      <= "111000000011010100001011100010101100011010001000111001100000101011001110110111010111101111001111101101110100011101101011000010010100110110110101010100";
reg_sig_51      <= "101011110101000010010000001110001111011110001000101100011100000010111100100111101110110101011100011111001100011110001010100101011100000001000111000100";
reg_sig_52      <= "111000101010110011010101010101111010110010000110011010011101010001100100110100000111110000111100111110001100111000111101001001001000011110001111010111";
reg_sig_53      <= "000001100100001111011010011000010101100111000111111110000111001001110110010110110010000011101001010101010101010110011101000100111110100110110011010010";
reg_sig_54      <= "100110000101000110110010011110100101110101011110100001110001111010110100111100000011110111101100110010000000100111010110110110010011000101111001110110";
reg_sig_55      <= "010101011101010101101111100000011111111001100010011001100001110110001011100010110000001111001110001110011000010100110001111111001101100001010010101111";
reg_sig_56      <= "000010000100110100000011000011001110110100011100010100100111001011010010100001101000010011100001001101101011011010111110100010111011011110101010010011";
reg_sig_57      <= "001011010100110000111100001111010010110101101101010100101011101010010001100001011111100000110010000111010111101111100110100100011010101010101010100101";
reg_sig_58      <= "010001111010101011110000100000011101001101110110111111110000000001101111000011000100101001001110010101111000001111000001100011010010101010011000001010";
reg_sig_59      <= "000011110110001000100011101101100111101100011010110010011010010000100010101011011001100000111001101010110011011111010111111111110011110001011110001011";
reg_sig_60      <= "110111110101011111110000100110010000010011111011100101111011111111001100100101011101100100000001000110010010100011100011110110010011100001000011011010";
reg_sig_61      <= "101010110010001010110011101011011001000111010100011110001011111111110000111001110100011010010100011001110100000010001100001001000001010111011011111001";
reg_sig_62      <= "111011011110000001110000000010100001000111001011000011100010010111010001111000111001001100011000011100111011111000010000001010100001101010110001101101";
reg_sig_63      <= "010101100110000100110110101110110010000010100010001110001010100010111101100111111100011000110000111111011000100101111001010000010011010110111111100001";
reg_sig_64      <= "111000010001011010101001100111001111010101010001000011111111001010010000010111111001011001000000110010111111010111101100110011111100010010000110101001";
reg_sig_65      <= "101111000001110101100001110000001110110110111110101010010100111010110101101111100011101110111110111100111010001011111001000000110110010010000100100011";
reg_sig_66      <= "011110001011110100110110101111011001111011100001100111001100100010110111001000011100101001000100111000111010100101110010100111100110001010000010111001";
reg_sig_67      <= "110110100001100011000111110011010111000110100011000101101101011101010011100010000011000001011010100010110011010110001100100101010111001000000101110110";
reg_sig_68      <= "100001010110100100010001001100101010001101010100001001100011001011000010010111101101100111010110010101000000100110011100101100001100001100110111000111";
reg_sig_69      <= "001011000110001111000110001011100001000101100111101110001000011101001001111100011100100100110010110001100010001100100001001111101110100110010001001001";
reg_sig_70      <= "101011101111100010000101000001010111101001010110100100111101010001010010100001100111111100111110001011100101111110100001001100011101111111011110101011";
reg_sig_71      <= "111011100011110101011001101000110000010110010000001011010111000011000100001000101010101001010001011000100010110110010011010111101111101000010100101011";
reg_sig_72      <= "101100001011101000001100000110100000100000111011011011100101100100011000010101001110100011000101000011001001010101111011001111111000000110101101010001";
reg_sig_73      <= "000010010000110011010111000111111111010111100001010111110100011100001111001111000110010001111001111010010110110001001011010010001000001100101000111100";
reg_sig_74      <= "101101010110111101000111011110111000111010100110010011010010010111011000100000101101011010100000110010101001100101110010001011110001010000111000100100";
reg_sig_75      <= "011100111010010101011000010111100101100011011100010000011010110110111010001100101101110110101100101001110100101111111101011110110100000010010010111110";
reg_sig_76      <= "010000100010111011101001101010100000000110011111000111100010110011001111101000111111001110011101010110110011001101100011000100100101000111011101011101";
reg_sig_77      <= "101000111100000111011100100011101110101110001110101011001110111000001011110100011101011101001111001100110111000111100100011101100001110000110000001001";
reg_sig_78      <= "000010011001100001110101110110001001100000000110000111011101111001000000100111000010110010000111011000101010111001110011111110010111001110010010100011";
reg_sig_79      <= "110101011111011101111011110001000111110000111000010110001011101100101101001110001011010010111011111010111100101010110101010110010100110101110001101011";
reg_sig_80      <= "101110101111000010010100000100111001100010111010110111001110001111101100000100100100010101101001100001011001000000101111110011110101001000110010010011";
reg_sig_81      <= "110101000101011100010001101110001110101001111010110100010011011010101001101110110110101010110000111100111111101100110000100001101011100110101101101011";
reg_sig_82      <= "011011011110001000010111010011111001001101010010000111011110011111001000001001000110111000011111010000010110010011011110010111000000110110010111111101";
reg_sig_83      <= "101111000110101111010011101101000111000100111110100000010111101000011010011101101100110101010101001011001101100001110010100111011001100111101100101101";
reg_sig_84      <= "001001000001000111111101000000000110100111100100000101111100110001110111010011110011000100000000110000000101100100111111101011111001111100110010100101";
reg_sig_85      <= "000011011111001010101111101000111010000100110000110101101001011101010011011101101010110000100100101100010111011110111011001011001110100101101111100110";
reg_sig_86      <= "011100011011000001010010111110010010101101011010010101011100101000011111010000101001110111011100100101110000101111000111110100110101010101111101101011";
reg_sig_87      <= "010100011101101001001110100010111101011100101100110001010011100101010100001101100110000011100010001111010010100101111000010011011010000011000011000011";
reg_sig_88      <= "101110100010010011110011010000100110000101110000110001110111011111110100111011111111101000001110010011010111110010100101100101101100001100010001111110";
reg_sig_89      <= "011010110100110011100110000111000101101100110011000110010000101000111101100001000111110000110110111110010101100010110000000101100100000110111001101111";
reg_sig_90      <= "101011000010000101011110000001010100101101101100111011100011000110010001010010010001110011001000001110110011000000100001110101011110000100010000010101";
reg_sig_91      <= "001010101001010111110101010000101010000010011100000101000010001010101010011010100100011001100001011110100111101010001111101010011110010111111110100110";
reg_sig_92      <= "010010111010110110110111101001011010110010101001010010111100110011000011101000101010101001010010111100110101111010010001111111101000011001110110001100";
reg_sig_93      <= "100000011100011010101010000011010111101110111100011011101100011101011010011110100101010000110101100001101111100111110110011100000101101001111000101011";
reg_sig_94      <= "010000010000010000011000100000000011101101111001110000111011110110000110101111101010100111011010011001001011110101101100001111110010001011011111100001";
reg_sig_95      <= "100011110110011001000000101100110010001010011011100010101001001001011011101010010111100011001100100010001111101001100001001010011100111010000111111101";
reg_sig_96      <= "000001101001111010101000111111001100111001000101001001110101001011010101010101000001110000011010011110000011100110010011111100100111010010010001100100";
reg_sig_97      <= "001000001111110101010100110011011011101100111000000000010000101001101010000000011001010010010111010000011001101101100011100010000111110011100111001001";
reg_sig_98      <= "101100011111001110010011011010000001110101000001100001011010000001100010100001101011010110010010100101111010110101000110011100111011110110010100111001";
reg_sig_99      <= "101110001111100011001000001101000001111001100100110011101110011010110111000010111011011111111011011001101011001111011111111010111001101100101001110011";

		elsif start= '1' then	
		codeword_avail <= '1';	
		end if;
	end if;
end process;
end rtl;